* Lumped Transmission Line Model
* Length: 0.6925m, Segments: 37549
* L/segment: 1.156e-11H, C/segment: 7.858e-16F

.param L_segment=1.1558457727310058e-11
.param C_segment=7.858283209454848e-16

.include Segment.sub

* Instantiation 37549 segments
X0 Vin N1 Segment
X1 N1 N2 Segment
X2 N2 N3 Segment
X3 N3 N4 Segment
X4 N4 N5 Segment
X5 N5 N6 Segment
X6 N6 N7 Segment
X7 N7 N8 Segment
X8 N8 N9 Segment
X9 N9 N10 Segment
X10 N10 N11 Segment
X11 N11 N12 Segment
X12 N12 N13 Segment
X13 N13 N14 Segment
X14 N14 N15 Segment
X15 N15 N16 Segment
X16 N16 N17 Segment
X17 N17 N18 Segment
X18 N18 N19 Segment
X19 N19 N20 Segment
X20 N20 N21 Segment
X21 N21 N22 Segment
X22 N22 N23 Segment
X23 N23 N24 Segment
X24 N24 N25 Segment
X25 N25 N26 Segment
X26 N26 N27 Segment
X27 N27 N28 Segment
X28 N28 N29 Segment
X29 N29 N30 Segment
X30 N30 N31 Segment
X31 N31 N32 Segment
X32 N32 N33 Segment
X33 N33 N34 Segment
X34 N34 N35 Segment
X35 N35 N36 Segment
X36 N36 N37 Segment
X37 N37 N38 Segment
X38 N38 N39 Segment
X39 N39 N40 Segment
X40 N40 N41 Segment
X41 N41 N42 Segment
X42 N42 N43 Segment
X43 N43 N44 Segment
X44 N44 N45 Segment
X45 N45 N46 Segment
X46 N46 N47 Segment
X47 N47 N48 Segment
X48 N48 N49 Segment
X49 N49 N50 Segment
X50 N50 N51 Segment
X51 N51 N52 Segment
X52 N52 N53 Segment
X53 N53 N54 Segment
X54 N54 N55 Segment
X55 N55 N56 Segment
X56 N56 N57 Segment
X57 N57 N58 Segment
X58 N58 N59 Segment
X59 N59 N60 Segment
X60 N60 N61 Segment
X61 N61 N62 Segment
X62 N62 N63 Segment
X63 N63 N64 Segment
X64 N64 N65 Segment
X65 N65 N66 Segment
X66 N66 N67 Segment
X67 N67 N68 Segment
X68 N68 N69 Segment
X69 N69 N70 Segment
X70 N70 N71 Segment
X71 N71 N72 Segment
X72 N72 N73 Segment
X73 N73 N74 Segment
X74 N74 N75 Segment
X75 N75 N76 Segment
X76 N76 N77 Segment
X77 N77 N78 Segment
X78 N78 N79 Segment
X79 N79 N80 Segment
X80 N80 N81 Segment
X81 N81 N82 Segment
X82 N82 N83 Segment
X83 N83 N84 Segment
X84 N84 N85 Segment
X85 N85 N86 Segment
X86 N86 N87 Segment
X87 N87 N88 Segment
X88 N88 N89 Segment
X89 N89 N90 Segment
X90 N90 N91 Segment
X91 N91 N92 Segment
X92 N92 N93 Segment
X93 N93 N94 Segment
X94 N94 N95 Segment
X95 N95 N96 Segment
X96 N96 N97 Segment
X97 N97 N98 Segment
X98 N98 N99 Segment
X99 N99 N100 Segment
X100 N100 N101 Segment
X101 N101 N102 Segment
X102 N102 N103 Segment
X103 N103 N104 Segment
X104 N104 N105 Segment
X105 N105 N106 Segment
X106 N106 N107 Segment
X107 N107 N108 Segment
X108 N108 N109 Segment
X109 N109 N110 Segment
X110 N110 N111 Segment
X111 N111 N112 Segment
X112 N112 N113 Segment
X113 N113 N114 Segment
X114 N114 N115 Segment
X115 N115 N116 Segment
X116 N116 N117 Segment
X117 N117 N118 Segment
X118 N118 N119 Segment
X119 N119 N120 Segment
X120 N120 N121 Segment
X121 N121 N122 Segment
X122 N122 N123 Segment
X123 N123 N124 Segment
X124 N124 N125 Segment
X125 N125 N126 Segment
X126 N126 N127 Segment
X127 N127 N128 Segment
X128 N128 N129 Segment
X129 N129 N130 Segment
X130 N130 N131 Segment
X131 N131 N132 Segment
X132 N132 N133 Segment
X133 N133 N134 Segment
X134 N134 N135 Segment
X135 N135 N136 Segment
X136 N136 N137 Segment
X137 N137 N138 Segment
X138 N138 N139 Segment
X139 N139 N140 Segment
X140 N140 N141 Segment
X141 N141 N142 Segment
X142 N142 N143 Segment
X143 N143 N144 Segment
X144 N144 N145 Segment
X145 N145 N146 Segment
X146 N146 N147 Segment
X147 N147 N148 Segment
X148 N148 N149 Segment
X149 N149 N150 Segment
X150 N150 N151 Segment
X151 N151 N152 Segment
X152 N152 N153 Segment
X153 N153 N154 Segment
X154 N154 N155 Segment
X155 N155 N156 Segment
X156 N156 N157 Segment
X157 N157 N158 Segment
X158 N158 N159 Segment
X159 N159 N160 Segment
X160 N160 N161 Segment
X161 N161 N162 Segment
X162 N162 N163 Segment
X163 N163 N164 Segment
X164 N164 N165 Segment
X165 N165 N166 Segment
X166 N166 N167 Segment
X167 N167 N168 Segment
X168 N168 N169 Segment
X169 N169 N170 Segment
X170 N170 N171 Segment
X171 N171 N172 Segment
X172 N172 N173 Segment
X173 N173 N174 Segment
X174 N174 N175 Segment
X175 N175 N176 Segment
X176 N176 N177 Segment
X177 N177 N178 Segment
X178 N178 N179 Segment
X179 N179 N180 Segment
X180 N180 N181 Segment
X181 N181 N182 Segment
X182 N182 N183 Segment
X183 N183 N184 Segment
X184 N184 N185 Segment
X185 N185 N186 Segment
X186 N186 N187 Segment
X187 N187 N188 Segment
X188 N188 N189 Segment
X189 N189 N190 Segment
X190 N190 N191 Segment
X191 N191 N192 Segment
X192 N192 N193 Segment
X193 N193 N194 Segment
X194 N194 N195 Segment
X195 N195 N196 Segment
X196 N196 N197 Segment
X197 N197 N198 Segment
X198 N198 N199 Segment
X199 N199 N200 Segment
X200 N200 N201 Segment
X201 N201 N202 Segment
X202 N202 N203 Segment
X203 N203 N204 Segment
X204 N204 N205 Segment
X205 N205 N206 Segment
X206 N206 N207 Segment
X207 N207 N208 Segment
X208 N208 N209 Segment
X209 N209 N210 Segment
X210 N210 N211 Segment
X211 N211 N212 Segment
X212 N212 N213 Segment
X213 N213 N214 Segment
X214 N214 N215 Segment
X215 N215 N216 Segment
X216 N216 N217 Segment
X217 N217 N218 Segment
X218 N218 N219 Segment
X219 N219 N220 Segment
X220 N220 N221 Segment
X221 N221 N222 Segment
X222 N222 N223 Segment
X223 N223 N224 Segment
X224 N224 N225 Segment
X225 N225 N226 Segment
X226 N226 N227 Segment
X227 N227 N228 Segment
X228 N228 N229 Segment
X229 N229 N230 Segment
X230 N230 N231 Segment
X231 N231 N232 Segment
X232 N232 N233 Segment
X233 N233 N234 Segment
X234 N234 N235 Segment
X235 N235 N236 Segment
X236 N236 N237 Segment
X237 N237 N238 Segment
X238 N238 N239 Segment
X239 N239 N240 Segment
X240 N240 N241 Segment
X241 N241 N242 Segment
X242 N242 N243 Segment
X243 N243 N244 Segment
X244 N244 N245 Segment
X245 N245 N246 Segment
X246 N246 N247 Segment
X247 N247 N248 Segment
X248 N248 N249 Segment
X249 N249 N250 Segment
X250 N250 N251 Segment
X251 N251 N252 Segment
X252 N252 N253 Segment
X253 N253 N254 Segment
X254 N254 N255 Segment
X255 N255 N256 Segment
X256 N256 N257 Segment
X257 N257 N258 Segment
X258 N258 N259 Segment
X259 N259 N260 Segment
X260 N260 N261 Segment
X261 N261 N262 Segment
X262 N262 N263 Segment
X263 N263 N264 Segment
X264 N264 N265 Segment
X265 N265 N266 Segment
X266 N266 N267 Segment
X267 N267 N268 Segment
X268 N268 N269 Segment
X269 N269 N270 Segment
X270 N270 N271 Segment
X271 N271 N272 Segment
X272 N272 N273 Segment
X273 N273 N274 Segment
X274 N274 N275 Segment
X275 N275 N276 Segment
X276 N276 N277 Segment
X277 N277 N278 Segment
X278 N278 N279 Segment
X279 N279 N280 Segment
X280 N280 N281 Segment
X281 N281 N282 Segment
X282 N282 N283 Segment
X283 N283 N284 Segment
X284 N284 N285 Segment
X285 N285 N286 Segment
X286 N286 N287 Segment
X287 N287 N288 Segment
X288 N288 N289 Segment
X289 N289 N290 Segment
X290 N290 N291 Segment
X291 N291 N292 Segment
X292 N292 N293 Segment
X293 N293 N294 Segment
X294 N294 N295 Segment
X295 N295 N296 Segment
X296 N296 N297 Segment
X297 N297 N298 Segment
X298 N298 N299 Segment
X299 N299 N300 Segment
X300 N300 N301 Segment
X301 N301 N302 Segment
X302 N302 N303 Segment
X303 N303 N304 Segment
X304 N304 N305 Segment
X305 N305 N306 Segment
X306 N306 N307 Segment
X307 N307 N308 Segment
X308 N308 N309 Segment
X309 N309 N310 Segment
X310 N310 N311 Segment
X311 N311 N312 Segment
X312 N312 N313 Segment
X313 N313 N314 Segment
X314 N314 N315 Segment
X315 N315 N316 Segment
X316 N316 N317 Segment
X317 N317 N318 Segment
X318 N318 N319 Segment
X319 N319 N320 Segment
X320 N320 N321 Segment
X321 N321 N322 Segment
X322 N322 N323 Segment
X323 N323 N324 Segment
X324 N324 N325 Segment
X325 N325 N326 Segment
X326 N326 N327 Segment
X327 N327 N328 Segment
X328 N328 N329 Segment
X329 N329 N330 Segment
X330 N330 N331 Segment
X331 N331 N332 Segment
X332 N332 N333 Segment
X333 N333 N334 Segment
X334 N334 N335 Segment
X335 N335 N336 Segment
X336 N336 N337 Segment
X337 N337 N338 Segment
X338 N338 N339 Segment
X339 N339 N340 Segment
X340 N340 N341 Segment
X341 N341 N342 Segment
X342 N342 N343 Segment
X343 N343 N344 Segment
X344 N344 N345 Segment
X345 N345 N346 Segment
X346 N346 N347 Segment
X347 N347 N348 Segment
X348 N348 N349 Segment
X349 N349 N350 Segment
X350 N350 N351 Segment
X351 N351 N352 Segment
X352 N352 N353 Segment
X353 N353 N354 Segment
X354 N354 N355 Segment
X355 N355 N356 Segment
X356 N356 N357 Segment
X357 N357 N358 Segment
X358 N358 N359 Segment
X359 N359 N360 Segment
X360 N360 N361 Segment
X361 N361 N362 Segment
X362 N362 N363 Segment
X363 N363 N364 Segment
X364 N364 N365 Segment
X365 N365 N366 Segment
X366 N366 N367 Segment
X367 N367 N368 Segment
X368 N368 N369 Segment
X369 N369 N370 Segment
X370 N370 N371 Segment
X371 N371 N372 Segment
X372 N372 N373 Segment
X373 N373 N374 Segment
X374 N374 N375 Segment
X375 N375 N376 Segment
X376 N376 N377 Segment
X377 N377 N378 Segment
X378 N378 N379 Segment
X379 N379 N380 Segment
X380 N380 N381 Segment
X381 N381 N382 Segment
X382 N382 N383 Segment
X383 N383 N384 Segment
X384 N384 N385 Segment
X385 N385 N386 Segment
X386 N386 N387 Segment
X387 N387 N388 Segment
X388 N388 N389 Segment
X389 N389 N390 Segment
X390 N390 N391 Segment
X391 N391 N392 Segment
X392 N392 N393 Segment
X393 N393 N394 Segment
X394 N394 N395 Segment
X395 N395 N396 Segment
X396 N396 N397 Segment
X397 N397 N398 Segment
X398 N398 N399 Segment
X399 N399 N400 Segment
X400 N400 N401 Segment
X401 N401 N402 Segment
X402 N402 N403 Segment
X403 N403 N404 Segment
X404 N404 N405 Segment
X405 N405 N406 Segment
X406 N406 N407 Segment
X407 N407 N408 Segment
X408 N408 N409 Segment
X409 N409 N410 Segment
X410 N410 N411 Segment
X411 N411 N412 Segment
X412 N412 N413 Segment
X413 N413 N414 Segment
X414 N414 N415 Segment
X415 N415 N416 Segment
X416 N416 N417 Segment
X417 N417 N418 Segment
X418 N418 N419 Segment
X419 N419 N420 Segment
X420 N420 N421 Segment
X421 N421 N422 Segment
X422 N422 N423 Segment
X423 N423 N424 Segment
X424 N424 N425 Segment
X425 N425 N426 Segment
X426 N426 N427 Segment
X427 N427 N428 Segment
X428 N428 N429 Segment
X429 N429 N430 Segment
X430 N430 N431 Segment
X431 N431 N432 Segment
X432 N432 N433 Segment
X433 N433 N434 Segment
X434 N434 N435 Segment
X435 N435 N436 Segment
X436 N436 N437 Segment
X437 N437 N438 Segment
X438 N438 N439 Segment
X439 N439 N440 Segment
X440 N440 N441 Segment
X441 N441 N442 Segment
X442 N442 N443 Segment
X443 N443 N444 Segment
X444 N444 N445 Segment
X445 N445 N446 Segment
X446 N446 N447 Segment
X447 N447 N448 Segment
X448 N448 N449 Segment
X449 N449 N450 Segment
X450 N450 N451 Segment
X451 N451 N452 Segment
X452 N452 N453 Segment
X453 N453 N454 Segment
X454 N454 N455 Segment
X455 N455 N456 Segment
X456 N456 N457 Segment
X457 N457 N458 Segment
X458 N458 N459 Segment
X459 N459 N460 Segment
X460 N460 N461 Segment
X461 N461 N462 Segment
X462 N462 N463 Segment
X463 N463 N464 Segment
X464 N464 N465 Segment
X465 N465 N466 Segment
X466 N466 N467 Segment
X467 N467 N468 Segment
X468 N468 N469 Segment
X469 N469 N470 Segment
X470 N470 N471 Segment
X471 N471 N472 Segment
X472 N472 N473 Segment
X473 N473 N474 Segment
X474 N474 N475 Segment
X475 N475 N476 Segment
X476 N476 N477 Segment
X477 N477 N478 Segment
X478 N478 N479 Segment
X479 N479 N480 Segment
X480 N480 N481 Segment
X481 N481 N482 Segment
X482 N482 N483 Segment
X483 N483 N484 Segment
X484 N484 N485 Segment
X485 N485 N486 Segment
X486 N486 N487 Segment
X487 N487 N488 Segment
X488 N488 N489 Segment
X489 N489 N490 Segment
X490 N490 N491 Segment
X491 N491 N492 Segment
X492 N492 N493 Segment
X493 N493 N494 Segment
X494 N494 N495 Segment
X495 N495 N496 Segment
X496 N496 N497 Segment
X497 N497 N498 Segment
X498 N498 N499 Segment
X499 N499 N500 Segment
X500 N500 N501 Segment
X501 N501 N502 Segment
X502 N502 N503 Segment
X503 N503 N504 Segment
X504 N504 N505 Segment
X505 N505 N506 Segment
X506 N506 N507 Segment
X507 N507 N508 Segment
X508 N508 N509 Segment
X509 N509 N510 Segment
X510 N510 N511 Segment
X511 N511 N512 Segment
X512 N512 N513 Segment
X513 N513 N514 Segment
X514 N514 N515 Segment
X515 N515 N516 Segment
X516 N516 N517 Segment
X517 N517 N518 Segment
X518 N518 N519 Segment
X519 N519 N520 Segment
X520 N520 N521 Segment
X521 N521 N522 Segment
X522 N522 N523 Segment
X523 N523 N524 Segment
X524 N524 N525 Segment
X525 N525 N526 Segment
X526 N526 N527 Segment
X527 N527 N528 Segment
X528 N528 N529 Segment
X529 N529 N530 Segment
X530 N530 N531 Segment
X531 N531 N532 Segment
X532 N532 N533 Segment
X533 N533 N534 Segment
X534 N534 N535 Segment
X535 N535 N536 Segment
X536 N536 N537 Segment
X537 N537 N538 Segment
X538 N538 N539 Segment
X539 N539 N540 Segment
X540 N540 N541 Segment
X541 N541 N542 Segment
X542 N542 N543 Segment
X543 N543 N544 Segment
X544 N544 N545 Segment
X545 N545 N546 Segment
X546 N546 N547 Segment
X547 N547 N548 Segment
X548 N548 N549 Segment
X549 N549 N550 Segment
X550 N550 N551 Segment
X551 N551 N552 Segment
X552 N552 N553 Segment
X553 N553 N554 Segment
X554 N554 N555 Segment
X555 N555 N556 Segment
X556 N556 N557 Segment
X557 N557 N558 Segment
X558 N558 N559 Segment
X559 N559 N560 Segment
X560 N560 N561 Segment
X561 N561 N562 Segment
X562 N562 N563 Segment
X563 N563 N564 Segment
X564 N564 N565 Segment
X565 N565 N566 Segment
X566 N566 N567 Segment
X567 N567 N568 Segment
X568 N568 N569 Segment
X569 N569 N570 Segment
X570 N570 N571 Segment
X571 N571 N572 Segment
X572 N572 N573 Segment
X573 N573 N574 Segment
X574 N574 N575 Segment
X575 N575 N576 Segment
X576 N576 N577 Segment
X577 N577 N578 Segment
X578 N578 N579 Segment
X579 N579 N580 Segment
X580 N580 N581 Segment
X581 N581 N582 Segment
X582 N582 N583 Segment
X583 N583 N584 Segment
X584 N584 N585 Segment
X585 N585 N586 Segment
X586 N586 N587 Segment
X587 N587 N588 Segment
X588 N588 N589 Segment
X589 N589 N590 Segment
X590 N590 N591 Segment
X591 N591 N592 Segment
X592 N592 N593 Segment
X593 N593 N594 Segment
X594 N594 N595 Segment
X595 N595 N596 Segment
X596 N596 N597 Segment
X597 N597 N598 Segment
X598 N598 N599 Segment
X599 N599 N600 Segment
X600 N600 N601 Segment
X601 N601 N602 Segment
X602 N602 N603 Segment
X603 N603 N604 Segment
X604 N604 N605 Segment
X605 N605 N606 Segment
X606 N606 N607 Segment
X607 N607 N608 Segment
X608 N608 N609 Segment
X609 N609 N610 Segment
X610 N610 N611 Segment
X611 N611 N612 Segment
X612 N612 N613 Segment
X613 N613 N614 Segment
X614 N614 N615 Segment
X615 N615 N616 Segment
X616 N616 N617 Segment
X617 N617 N618 Segment
X618 N618 N619 Segment
X619 N619 N620 Segment
X620 N620 N621 Segment
X621 N621 N622 Segment
X622 N622 N623 Segment
X623 N623 N624 Segment
X624 N624 N625 Segment
X625 N625 N626 Segment
X626 N626 N627 Segment
X627 N627 N628 Segment
X628 N628 N629 Segment
X629 N629 N630 Segment
X630 N630 N631 Segment
X631 N631 N632 Segment
X632 N632 N633 Segment
X633 N633 N634 Segment
X634 N634 N635 Segment
X635 N635 N636 Segment
X636 N636 N637 Segment
X637 N637 N638 Segment
X638 N638 N639 Segment
X639 N639 N640 Segment
X640 N640 N641 Segment
X641 N641 N642 Segment
X642 N642 N643 Segment
X643 N643 N644 Segment
X644 N644 N645 Segment
X645 N645 N646 Segment
X646 N646 N647 Segment
X647 N647 N648 Segment
X648 N648 N649 Segment
X649 N649 N650 Segment
X650 N650 N651 Segment
X651 N651 N652 Segment
X652 N652 N653 Segment
X653 N653 N654 Segment
X654 N654 N655 Segment
X655 N655 N656 Segment
X656 N656 N657 Segment
X657 N657 N658 Segment
X658 N658 N659 Segment
X659 N659 N660 Segment
X660 N660 N661 Segment
X661 N661 N662 Segment
X662 N662 N663 Segment
X663 N663 N664 Segment
X664 N664 N665 Segment
X665 N665 N666 Segment
X666 N666 N667 Segment
X667 N667 N668 Segment
X668 N668 N669 Segment
X669 N669 N670 Segment
X670 N670 N671 Segment
X671 N671 N672 Segment
X672 N672 N673 Segment
X673 N673 N674 Segment
X674 N674 N675 Segment
X675 N675 N676 Segment
X676 N676 N677 Segment
X677 N677 N678 Segment
X678 N678 N679 Segment
X679 N679 N680 Segment
X680 N680 N681 Segment
X681 N681 N682 Segment
X682 N682 N683 Segment
X683 N683 N684 Segment
X684 N684 N685 Segment
X685 N685 N686 Segment
X686 N686 N687 Segment
X687 N687 N688 Segment
X688 N688 N689 Segment
X689 N689 N690 Segment
X690 N690 N691 Segment
X691 N691 N692 Segment
X692 N692 N693 Segment
X693 N693 N694 Segment
X694 N694 N695 Segment
X695 N695 N696 Segment
X696 N696 N697 Segment
X697 N697 N698 Segment
X698 N698 N699 Segment
X699 N699 N700 Segment
X700 N700 N701 Segment
X701 N701 N702 Segment
X702 N702 N703 Segment
X703 N703 N704 Segment
X704 N704 N705 Segment
X705 N705 N706 Segment
X706 N706 N707 Segment
X707 N707 N708 Segment
X708 N708 N709 Segment
X709 N709 N710 Segment
X710 N710 N711 Segment
X711 N711 N712 Segment
X712 N712 N713 Segment
X713 N713 N714 Segment
X714 N714 N715 Segment
X715 N715 N716 Segment
X716 N716 N717 Segment
X717 N717 N718 Segment
X718 N718 N719 Segment
X719 N719 N720 Segment
X720 N720 N721 Segment
X721 N721 N722 Segment
X722 N722 N723 Segment
X723 N723 N724 Segment
X724 N724 N725 Segment
X725 N725 N726 Segment
X726 N726 N727 Segment
X727 N727 N728 Segment
X728 N728 N729 Segment
X729 N729 N730 Segment
X730 N730 N731 Segment
X731 N731 N732 Segment
X732 N732 N733 Segment
X733 N733 N734 Segment
X734 N734 N735 Segment
X735 N735 N736 Segment
X736 N736 N737 Segment
X737 N737 N738 Segment
X738 N738 N739 Segment
X739 N739 N740 Segment
X740 N740 N741 Segment
X741 N741 N742 Segment
X742 N742 N743 Segment
X743 N743 N744 Segment
X744 N744 N745 Segment
X745 N745 N746 Segment
X746 N746 N747 Segment
X747 N747 N748 Segment
X748 N748 N749 Segment
X749 N749 N750 Segment
X750 N750 N751 Segment
X751 N751 N752 Segment
X752 N752 N753 Segment
X753 N753 N754 Segment
X754 N754 N755 Segment
X755 N755 N756 Segment
X756 N756 N757 Segment
X757 N757 N758 Segment
X758 N758 N759 Segment
X759 N759 N760 Segment
X760 N760 N761 Segment
X761 N761 N762 Segment
X762 N762 N763 Segment
X763 N763 N764 Segment
X764 N764 N765 Segment
X765 N765 N766 Segment
X766 N766 N767 Segment
X767 N767 N768 Segment
X768 N768 N769 Segment
X769 N769 N770 Segment
X770 N770 N771 Segment
X771 N771 N772 Segment
X772 N772 N773 Segment
X773 N773 N774 Segment
X774 N774 N775 Segment
X775 N775 N776 Segment
X776 N776 N777 Segment
X777 N777 N778 Segment
X778 N778 N779 Segment
X779 N779 N780 Segment
X780 N780 N781 Segment
X781 N781 N782 Segment
X782 N782 N783 Segment
X783 N783 N784 Segment
X784 N784 N785 Segment
X785 N785 N786 Segment
X786 N786 N787 Segment
X787 N787 N788 Segment
X788 N788 N789 Segment
X789 N789 N790 Segment
X790 N790 N791 Segment
X791 N791 N792 Segment
X792 N792 N793 Segment
X793 N793 N794 Segment
X794 N794 N795 Segment
X795 N795 N796 Segment
X796 N796 N797 Segment
X797 N797 N798 Segment
X798 N798 N799 Segment
X799 N799 N800 Segment
X800 N800 N801 Segment
X801 N801 N802 Segment
X802 N802 N803 Segment
X803 N803 N804 Segment
X804 N804 N805 Segment
X805 N805 N806 Segment
X806 N806 N807 Segment
X807 N807 N808 Segment
X808 N808 N809 Segment
X809 N809 N810 Segment
X810 N810 N811 Segment
X811 N811 N812 Segment
X812 N812 N813 Segment
X813 N813 N814 Segment
X814 N814 N815 Segment
X815 N815 N816 Segment
X816 N816 N817 Segment
X817 N817 N818 Segment
X818 N818 N819 Segment
X819 N819 N820 Segment
X820 N820 N821 Segment
X821 N821 N822 Segment
X822 N822 N823 Segment
X823 N823 N824 Segment
X824 N824 N825 Segment
X825 N825 N826 Segment
X826 N826 N827 Segment
X827 N827 N828 Segment
X828 N828 N829 Segment
X829 N829 N830 Segment
X830 N830 N831 Segment
X831 N831 N832 Segment
X832 N832 N833 Segment
X833 N833 N834 Segment
X834 N834 N835 Segment
X835 N835 N836 Segment
X836 N836 N837 Segment
X837 N837 N838 Segment
X838 N838 N839 Segment
X839 N839 N840 Segment
X840 N840 N841 Segment
X841 N841 N842 Segment
X842 N842 N843 Segment
X843 N843 N844 Segment
X844 N844 N845 Segment
X845 N845 N846 Segment
X846 N846 N847 Segment
X847 N847 N848 Segment
X848 N848 N849 Segment
X849 N849 N850 Segment
X850 N850 N851 Segment
X851 N851 N852 Segment
X852 N852 N853 Segment
X853 N853 N854 Segment
X854 N854 N855 Segment
X855 N855 N856 Segment
X856 N856 N857 Segment
X857 N857 N858 Segment
X858 N858 N859 Segment
X859 N859 N860 Segment
X860 N860 N861 Segment
X861 N861 N862 Segment
X862 N862 N863 Segment
X863 N863 N864 Segment
X864 N864 N865 Segment
X865 N865 N866 Segment
X866 N866 N867 Segment
X867 N867 N868 Segment
X868 N868 N869 Segment
X869 N869 N870 Segment
X870 N870 N871 Segment
X871 N871 N872 Segment
X872 N872 N873 Segment
X873 N873 N874 Segment
X874 N874 N875 Segment
X875 N875 N876 Segment
X876 N876 N877 Segment
X877 N877 N878 Segment
X878 N878 N879 Segment
X879 N879 N880 Segment
X880 N880 N881 Segment
X881 N881 N882 Segment
X882 N882 N883 Segment
X883 N883 N884 Segment
X884 N884 N885 Segment
X885 N885 N886 Segment
X886 N886 N887 Segment
X887 N887 N888 Segment
X888 N888 N889 Segment
X889 N889 N890 Segment
X890 N890 N891 Segment
X891 N891 N892 Segment
X892 N892 N893 Segment
X893 N893 N894 Segment
X894 N894 N895 Segment
X895 N895 N896 Segment
X896 N896 N897 Segment
X897 N897 N898 Segment
X898 N898 N899 Segment
X899 N899 N900 Segment
X900 N900 N901 Segment
X901 N901 N902 Segment
X902 N902 N903 Segment
X903 N903 N904 Segment
X904 N904 N905 Segment
X905 N905 N906 Segment
X906 N906 N907 Segment
X907 N907 N908 Segment
X908 N908 N909 Segment
X909 N909 N910 Segment
X910 N910 N911 Segment
X911 N911 N912 Segment
X912 N912 N913 Segment
X913 N913 N914 Segment
X914 N914 N915 Segment
X915 N915 N916 Segment
X916 N916 N917 Segment
X917 N917 N918 Segment
X918 N918 N919 Segment
X919 N919 N920 Segment
X920 N920 N921 Segment
X921 N921 N922 Segment
X922 N922 N923 Segment
X923 N923 N924 Segment
X924 N924 N925 Segment
X925 N925 N926 Segment
X926 N926 N927 Segment
X927 N927 N928 Segment
X928 N928 N929 Segment
X929 N929 N930 Segment
X930 N930 N931 Segment
X931 N931 N932 Segment
X932 N932 N933 Segment
X933 N933 N934 Segment
X934 N934 N935 Segment
X935 N935 N936 Segment
X936 N936 N937 Segment
X937 N937 N938 Segment
X938 N938 N939 Segment
X939 N939 N940 Segment
X940 N940 N941 Segment
X941 N941 N942 Segment
X942 N942 N943 Segment
X943 N943 N944 Segment
X944 N944 N945 Segment
X945 N945 N946 Segment
X946 N946 N947 Segment
X947 N947 N948 Segment
X948 N948 N949 Segment
X949 N949 N950 Segment
X950 N950 N951 Segment
X951 N951 N952 Segment
X952 N952 N953 Segment
X953 N953 N954 Segment
X954 N954 N955 Segment
X955 N955 N956 Segment
X956 N956 N957 Segment
X957 N957 N958 Segment
X958 N958 N959 Segment
X959 N959 N960 Segment
X960 N960 N961 Segment
X961 N961 N962 Segment
X962 N962 N963 Segment
X963 N963 N964 Segment
X964 N964 N965 Segment
X965 N965 N966 Segment
X966 N966 N967 Segment
X967 N967 N968 Segment
X968 N968 N969 Segment
X969 N969 N970 Segment
X970 N970 N971 Segment
X971 N971 N972 Segment
X972 N972 N973 Segment
X973 N973 N974 Segment
X974 N974 N975 Segment
X975 N975 N976 Segment
X976 N976 N977 Segment
X977 N977 N978 Segment
X978 N978 N979 Segment
X979 N979 N980 Segment
X980 N980 N981 Segment
X981 N981 N982 Segment
X982 N982 N983 Segment
X983 N983 N984 Segment
X984 N984 N985 Segment
X985 N985 N986 Segment
X986 N986 N987 Segment
X987 N987 N988 Segment
X988 N988 N989 Segment
X989 N989 N990 Segment
X990 N990 N991 Segment
X991 N991 N992 Segment
X992 N992 N993 Segment
X993 N993 N994 Segment
X994 N994 N995 Segment
X995 N995 N996 Segment
X996 N996 N997 Segment
X997 N997 N998 Segment
X998 N998 N999 Segment
X999 N999 N1000 Segment
X1000 N1000 N1001 Segment
X1001 N1001 N1002 Segment
X1002 N1002 N1003 Segment
X1003 N1003 N1004 Segment
X1004 N1004 N1005 Segment
X1005 N1005 N1006 Segment
X1006 N1006 N1007 Segment
X1007 N1007 N1008 Segment
X1008 N1008 N1009 Segment
X1009 N1009 N1010 Segment
X1010 N1010 N1011 Segment
X1011 N1011 N1012 Segment
X1012 N1012 N1013 Segment
X1013 N1013 N1014 Segment
X1014 N1014 N1015 Segment
X1015 N1015 N1016 Segment
X1016 N1016 N1017 Segment
X1017 N1017 N1018 Segment
X1018 N1018 N1019 Segment
X1019 N1019 N1020 Segment
X1020 N1020 N1021 Segment
X1021 N1021 N1022 Segment
X1022 N1022 N1023 Segment
X1023 N1023 N1024 Segment
X1024 N1024 N1025 Segment
X1025 N1025 N1026 Segment
X1026 N1026 N1027 Segment
X1027 N1027 N1028 Segment
X1028 N1028 N1029 Segment
X1029 N1029 N1030 Segment
X1030 N1030 N1031 Segment
X1031 N1031 N1032 Segment
X1032 N1032 N1033 Segment
X1033 N1033 N1034 Segment
X1034 N1034 N1035 Segment
X1035 N1035 N1036 Segment
X1036 N1036 N1037 Segment
X1037 N1037 N1038 Segment
X1038 N1038 N1039 Segment
X1039 N1039 N1040 Segment
X1040 N1040 N1041 Segment
X1041 N1041 N1042 Segment
X1042 N1042 N1043 Segment
X1043 N1043 N1044 Segment
X1044 N1044 N1045 Segment
X1045 N1045 N1046 Segment
X1046 N1046 N1047 Segment
X1047 N1047 N1048 Segment
X1048 N1048 N1049 Segment
X1049 N1049 N1050 Segment
X1050 N1050 N1051 Segment
X1051 N1051 N1052 Segment
X1052 N1052 N1053 Segment
X1053 N1053 N1054 Segment
X1054 N1054 N1055 Segment
X1055 N1055 N1056 Segment
X1056 N1056 N1057 Segment
X1057 N1057 N1058 Segment
X1058 N1058 N1059 Segment
X1059 N1059 N1060 Segment
X1060 N1060 N1061 Segment
X1061 N1061 N1062 Segment
X1062 N1062 N1063 Segment
X1063 N1063 N1064 Segment
X1064 N1064 N1065 Segment
X1065 N1065 N1066 Segment
X1066 N1066 N1067 Segment
X1067 N1067 N1068 Segment
X1068 N1068 N1069 Segment
X1069 N1069 N1070 Segment
X1070 N1070 N1071 Segment
X1071 N1071 N1072 Segment
X1072 N1072 N1073 Segment
X1073 N1073 N1074 Segment
X1074 N1074 N1075 Segment
X1075 N1075 N1076 Segment
X1076 N1076 N1077 Segment
X1077 N1077 N1078 Segment
X1078 N1078 N1079 Segment
X1079 N1079 N1080 Segment
X1080 N1080 N1081 Segment
X1081 N1081 N1082 Segment
X1082 N1082 N1083 Segment
X1083 N1083 N1084 Segment
X1084 N1084 N1085 Segment
X1085 N1085 N1086 Segment
X1086 N1086 N1087 Segment
X1087 N1087 N1088 Segment
X1088 N1088 N1089 Segment
X1089 N1089 N1090 Segment
X1090 N1090 N1091 Segment
X1091 N1091 N1092 Segment
X1092 N1092 N1093 Segment
X1093 N1093 N1094 Segment
X1094 N1094 N1095 Segment
X1095 N1095 N1096 Segment
X1096 N1096 N1097 Segment
X1097 N1097 N1098 Segment
X1098 N1098 N1099 Segment
X1099 N1099 N1100 Segment
X1100 N1100 N1101 Segment
X1101 N1101 N1102 Segment
X1102 N1102 N1103 Segment
X1103 N1103 N1104 Segment
X1104 N1104 N1105 Segment
X1105 N1105 N1106 Segment
X1106 N1106 N1107 Segment
X1107 N1107 N1108 Segment
X1108 N1108 N1109 Segment
X1109 N1109 N1110 Segment
X1110 N1110 N1111 Segment
X1111 N1111 N1112 Segment
X1112 N1112 N1113 Segment
X1113 N1113 N1114 Segment
X1114 N1114 N1115 Segment
X1115 N1115 N1116 Segment
X1116 N1116 N1117 Segment
X1117 N1117 N1118 Segment
X1118 N1118 N1119 Segment
X1119 N1119 N1120 Segment
X1120 N1120 N1121 Segment
X1121 N1121 N1122 Segment
X1122 N1122 N1123 Segment
X1123 N1123 N1124 Segment
X1124 N1124 N1125 Segment
X1125 N1125 N1126 Segment
X1126 N1126 N1127 Segment
X1127 N1127 N1128 Segment
X1128 N1128 N1129 Segment
X1129 N1129 N1130 Segment
X1130 N1130 N1131 Segment
X1131 N1131 N1132 Segment
X1132 N1132 N1133 Segment
X1133 N1133 N1134 Segment
X1134 N1134 N1135 Segment
X1135 N1135 N1136 Segment
X1136 N1136 N1137 Segment
X1137 N1137 N1138 Segment
X1138 N1138 N1139 Segment
X1139 N1139 N1140 Segment
X1140 N1140 N1141 Segment
X1141 N1141 N1142 Segment
X1142 N1142 N1143 Segment
X1143 N1143 N1144 Segment
X1144 N1144 N1145 Segment
X1145 N1145 N1146 Segment
X1146 N1146 N1147 Segment
X1147 N1147 N1148 Segment
X1148 N1148 N1149 Segment
X1149 N1149 N1150 Segment
X1150 N1150 N1151 Segment
X1151 N1151 N1152 Segment
X1152 N1152 N1153 Segment
X1153 N1153 N1154 Segment
X1154 N1154 N1155 Segment
X1155 N1155 N1156 Segment
X1156 N1156 N1157 Segment
X1157 N1157 N1158 Segment
X1158 N1158 N1159 Segment
X1159 N1159 N1160 Segment
X1160 N1160 N1161 Segment
X1161 N1161 N1162 Segment
X1162 N1162 N1163 Segment
X1163 N1163 N1164 Segment
X1164 N1164 N1165 Segment
X1165 N1165 N1166 Segment
X1166 N1166 N1167 Segment
X1167 N1167 N1168 Segment
X1168 N1168 N1169 Segment
X1169 N1169 N1170 Segment
X1170 N1170 N1171 Segment
X1171 N1171 N1172 Segment
X1172 N1172 N1173 Segment
X1173 N1173 N1174 Segment
X1174 N1174 N1175 Segment
X1175 N1175 N1176 Segment
X1176 N1176 N1177 Segment
X1177 N1177 N1178 Segment
X1178 N1178 N1179 Segment
X1179 N1179 N1180 Segment
X1180 N1180 N1181 Segment
X1181 N1181 N1182 Segment
X1182 N1182 N1183 Segment
X1183 N1183 N1184 Segment
X1184 N1184 N1185 Segment
X1185 N1185 N1186 Segment
X1186 N1186 N1187 Segment
X1187 N1187 N1188 Segment
X1188 N1188 N1189 Segment
X1189 N1189 N1190 Segment
X1190 N1190 N1191 Segment
X1191 N1191 N1192 Segment
X1192 N1192 N1193 Segment
X1193 N1193 N1194 Segment
X1194 N1194 N1195 Segment
X1195 N1195 N1196 Segment
X1196 N1196 N1197 Segment
X1197 N1197 N1198 Segment
X1198 N1198 N1199 Segment
X1199 N1199 N1200 Segment
X1200 N1200 N1201 Segment
X1201 N1201 N1202 Segment
X1202 N1202 N1203 Segment
X1203 N1203 N1204 Segment
X1204 N1204 N1205 Segment
X1205 N1205 N1206 Segment
X1206 N1206 N1207 Segment
X1207 N1207 N1208 Segment
X1208 N1208 N1209 Segment
X1209 N1209 N1210 Segment
X1210 N1210 N1211 Segment
X1211 N1211 N1212 Segment
X1212 N1212 N1213 Segment
X1213 N1213 N1214 Segment
X1214 N1214 N1215 Segment
X1215 N1215 N1216 Segment
X1216 N1216 N1217 Segment
X1217 N1217 N1218 Segment
X1218 N1218 N1219 Segment
X1219 N1219 N1220 Segment
X1220 N1220 N1221 Segment
X1221 N1221 N1222 Segment
X1222 N1222 N1223 Segment
X1223 N1223 N1224 Segment
X1224 N1224 N1225 Segment
X1225 N1225 N1226 Segment
X1226 N1226 N1227 Segment
X1227 N1227 N1228 Segment
X1228 N1228 N1229 Segment
X1229 N1229 N1230 Segment
X1230 N1230 N1231 Segment
X1231 N1231 N1232 Segment
X1232 N1232 N1233 Segment
X1233 N1233 N1234 Segment
X1234 N1234 N1235 Segment
X1235 N1235 N1236 Segment
X1236 N1236 N1237 Segment
X1237 N1237 N1238 Segment
X1238 N1238 N1239 Segment
X1239 N1239 N1240 Segment
X1240 N1240 N1241 Segment
X1241 N1241 N1242 Segment
X1242 N1242 N1243 Segment
X1243 N1243 N1244 Segment
X1244 N1244 N1245 Segment
X1245 N1245 N1246 Segment
X1246 N1246 N1247 Segment
X1247 N1247 N1248 Segment
X1248 N1248 N1249 Segment
X1249 N1249 N1250 Segment
X1250 N1250 N1251 Segment
X1251 N1251 N1252 Segment
X1252 N1252 N1253 Segment
X1253 N1253 N1254 Segment
X1254 N1254 N1255 Segment
X1255 N1255 N1256 Segment
X1256 N1256 N1257 Segment
X1257 N1257 N1258 Segment
X1258 N1258 N1259 Segment
X1259 N1259 N1260 Segment
X1260 N1260 N1261 Segment
X1261 N1261 N1262 Segment
X1262 N1262 N1263 Segment
X1263 N1263 N1264 Segment
X1264 N1264 N1265 Segment
X1265 N1265 N1266 Segment
X1266 N1266 N1267 Segment
X1267 N1267 N1268 Segment
X1268 N1268 N1269 Segment
X1269 N1269 N1270 Segment
X1270 N1270 N1271 Segment
X1271 N1271 N1272 Segment
X1272 N1272 N1273 Segment
X1273 N1273 N1274 Segment
X1274 N1274 N1275 Segment
X1275 N1275 N1276 Segment
X1276 N1276 N1277 Segment
X1277 N1277 N1278 Segment
X1278 N1278 N1279 Segment
X1279 N1279 N1280 Segment
X1280 N1280 N1281 Segment
X1281 N1281 N1282 Segment
X1282 N1282 N1283 Segment
X1283 N1283 N1284 Segment
X1284 N1284 N1285 Segment
X1285 N1285 N1286 Segment
X1286 N1286 N1287 Segment
X1287 N1287 N1288 Segment
X1288 N1288 N1289 Segment
X1289 N1289 N1290 Segment
X1290 N1290 N1291 Segment
X1291 N1291 N1292 Segment
X1292 N1292 N1293 Segment
X1293 N1293 N1294 Segment
X1294 N1294 N1295 Segment
X1295 N1295 N1296 Segment
X1296 N1296 N1297 Segment
X1297 N1297 N1298 Segment
X1298 N1298 N1299 Segment
X1299 N1299 N1300 Segment
X1300 N1300 N1301 Segment
X1301 N1301 N1302 Segment
X1302 N1302 N1303 Segment
X1303 N1303 N1304 Segment
X1304 N1304 N1305 Segment
X1305 N1305 N1306 Segment
X1306 N1306 N1307 Segment
X1307 N1307 N1308 Segment
X1308 N1308 N1309 Segment
X1309 N1309 N1310 Segment
X1310 N1310 N1311 Segment
X1311 N1311 N1312 Segment
X1312 N1312 N1313 Segment
X1313 N1313 N1314 Segment
X1314 N1314 N1315 Segment
X1315 N1315 N1316 Segment
X1316 N1316 N1317 Segment
X1317 N1317 N1318 Segment
X1318 N1318 N1319 Segment
X1319 N1319 N1320 Segment
X1320 N1320 N1321 Segment
X1321 N1321 N1322 Segment
X1322 N1322 N1323 Segment
X1323 N1323 N1324 Segment
X1324 N1324 N1325 Segment
X1325 N1325 N1326 Segment
X1326 N1326 N1327 Segment
X1327 N1327 N1328 Segment
X1328 N1328 N1329 Segment
X1329 N1329 N1330 Segment
X1330 N1330 N1331 Segment
X1331 N1331 N1332 Segment
X1332 N1332 N1333 Segment
X1333 N1333 N1334 Segment
X1334 N1334 N1335 Segment
X1335 N1335 N1336 Segment
X1336 N1336 N1337 Segment
X1337 N1337 N1338 Segment
X1338 N1338 N1339 Segment
X1339 N1339 N1340 Segment
X1340 N1340 N1341 Segment
X1341 N1341 N1342 Segment
X1342 N1342 N1343 Segment
X1343 N1343 N1344 Segment
X1344 N1344 N1345 Segment
X1345 N1345 N1346 Segment
X1346 N1346 N1347 Segment
X1347 N1347 N1348 Segment
X1348 N1348 N1349 Segment
X1349 N1349 N1350 Segment
X1350 N1350 N1351 Segment
X1351 N1351 N1352 Segment
X1352 N1352 N1353 Segment
X1353 N1353 N1354 Segment
X1354 N1354 N1355 Segment
X1355 N1355 N1356 Segment
X1356 N1356 N1357 Segment
X1357 N1357 N1358 Segment
X1358 N1358 N1359 Segment
X1359 N1359 N1360 Segment
X1360 N1360 N1361 Segment
X1361 N1361 N1362 Segment
X1362 N1362 N1363 Segment
X1363 N1363 N1364 Segment
X1364 N1364 N1365 Segment
X1365 N1365 N1366 Segment
X1366 N1366 N1367 Segment
X1367 N1367 N1368 Segment
X1368 N1368 N1369 Segment
X1369 N1369 N1370 Segment
X1370 N1370 N1371 Segment
X1371 N1371 N1372 Segment
X1372 N1372 N1373 Segment
X1373 N1373 N1374 Segment
X1374 N1374 N1375 Segment
X1375 N1375 N1376 Segment
X1376 N1376 N1377 Segment
X1377 N1377 N1378 Segment
X1378 N1378 N1379 Segment
X1379 N1379 N1380 Segment
X1380 N1380 N1381 Segment
X1381 N1381 N1382 Segment
X1382 N1382 N1383 Segment
X1383 N1383 N1384 Segment
X1384 N1384 N1385 Segment
X1385 N1385 N1386 Segment
X1386 N1386 N1387 Segment
X1387 N1387 N1388 Segment
X1388 N1388 N1389 Segment
X1389 N1389 N1390 Segment
X1390 N1390 N1391 Segment
X1391 N1391 N1392 Segment
X1392 N1392 N1393 Segment
X1393 N1393 N1394 Segment
X1394 N1394 N1395 Segment
X1395 N1395 N1396 Segment
X1396 N1396 N1397 Segment
X1397 N1397 N1398 Segment
X1398 N1398 N1399 Segment
X1399 N1399 N1400 Segment
X1400 N1400 N1401 Segment
X1401 N1401 N1402 Segment
X1402 N1402 N1403 Segment
X1403 N1403 N1404 Segment
X1404 N1404 N1405 Segment
X1405 N1405 N1406 Segment
X1406 N1406 N1407 Segment
X1407 N1407 N1408 Segment
X1408 N1408 N1409 Segment
X1409 N1409 N1410 Segment
X1410 N1410 N1411 Segment
X1411 N1411 N1412 Segment
X1412 N1412 N1413 Segment
X1413 N1413 N1414 Segment
X1414 N1414 N1415 Segment
X1415 N1415 N1416 Segment
X1416 N1416 N1417 Segment
X1417 N1417 N1418 Segment
X1418 N1418 N1419 Segment
X1419 N1419 N1420 Segment
X1420 N1420 N1421 Segment
X1421 N1421 N1422 Segment
X1422 N1422 N1423 Segment
X1423 N1423 N1424 Segment
X1424 N1424 N1425 Segment
X1425 N1425 N1426 Segment
X1426 N1426 N1427 Segment
X1427 N1427 N1428 Segment
X1428 N1428 N1429 Segment
X1429 N1429 N1430 Segment
X1430 N1430 N1431 Segment
X1431 N1431 N1432 Segment
X1432 N1432 N1433 Segment
X1433 N1433 N1434 Segment
X1434 N1434 N1435 Segment
X1435 N1435 N1436 Segment
X1436 N1436 N1437 Segment
X1437 N1437 N1438 Segment
X1438 N1438 N1439 Segment
X1439 N1439 N1440 Segment
X1440 N1440 N1441 Segment
X1441 N1441 N1442 Segment
X1442 N1442 N1443 Segment
X1443 N1443 N1444 Segment
X1444 N1444 N1445 Segment
X1445 N1445 N1446 Segment
X1446 N1446 N1447 Segment
X1447 N1447 N1448 Segment
X1448 N1448 N1449 Segment
X1449 N1449 N1450 Segment
X1450 N1450 N1451 Segment
X1451 N1451 N1452 Segment
X1452 N1452 N1453 Segment
X1453 N1453 N1454 Segment
X1454 N1454 N1455 Segment
X1455 N1455 N1456 Segment
X1456 N1456 N1457 Segment
X1457 N1457 N1458 Segment
X1458 N1458 N1459 Segment
X1459 N1459 N1460 Segment
X1460 N1460 N1461 Segment
X1461 N1461 N1462 Segment
X1462 N1462 N1463 Segment
X1463 N1463 N1464 Segment
X1464 N1464 N1465 Segment
X1465 N1465 N1466 Segment
X1466 N1466 N1467 Segment
X1467 N1467 N1468 Segment
X1468 N1468 N1469 Segment
X1469 N1469 N1470 Segment
X1470 N1470 N1471 Segment
X1471 N1471 N1472 Segment
X1472 N1472 N1473 Segment
X1473 N1473 N1474 Segment
X1474 N1474 N1475 Segment
X1475 N1475 N1476 Segment
X1476 N1476 N1477 Segment
X1477 N1477 N1478 Segment
X1478 N1478 N1479 Segment
X1479 N1479 N1480 Segment
X1480 N1480 N1481 Segment
X1481 N1481 N1482 Segment
X1482 N1482 N1483 Segment
X1483 N1483 N1484 Segment
X1484 N1484 N1485 Segment
X1485 N1485 N1486 Segment
X1486 N1486 N1487 Segment
X1487 N1487 N1488 Segment
X1488 N1488 N1489 Segment
X1489 N1489 N1490 Segment
X1490 N1490 N1491 Segment
X1491 N1491 N1492 Segment
X1492 N1492 N1493 Segment
X1493 N1493 N1494 Segment
X1494 N1494 N1495 Segment
X1495 N1495 N1496 Segment
X1496 N1496 N1497 Segment
X1497 N1497 N1498 Segment
X1498 N1498 N1499 Segment
X1499 N1499 N1500 Segment
X1500 N1500 N1501 Segment
X1501 N1501 N1502 Segment
X1502 N1502 N1503 Segment
X1503 N1503 N1504 Segment
X1504 N1504 N1505 Segment
X1505 N1505 N1506 Segment
X1506 N1506 N1507 Segment
X1507 N1507 N1508 Segment
X1508 N1508 N1509 Segment
X1509 N1509 N1510 Segment
X1510 N1510 N1511 Segment
X1511 N1511 N1512 Segment
X1512 N1512 N1513 Segment
X1513 N1513 N1514 Segment
X1514 N1514 N1515 Segment
X1515 N1515 N1516 Segment
X1516 N1516 N1517 Segment
X1517 N1517 N1518 Segment
X1518 N1518 N1519 Segment
X1519 N1519 N1520 Segment
X1520 N1520 N1521 Segment
X1521 N1521 N1522 Segment
X1522 N1522 N1523 Segment
X1523 N1523 N1524 Segment
X1524 N1524 N1525 Segment
X1525 N1525 N1526 Segment
X1526 N1526 N1527 Segment
X1527 N1527 N1528 Segment
X1528 N1528 N1529 Segment
X1529 N1529 N1530 Segment
X1530 N1530 N1531 Segment
X1531 N1531 N1532 Segment
X1532 N1532 N1533 Segment
X1533 N1533 N1534 Segment
X1534 N1534 N1535 Segment
X1535 N1535 N1536 Segment
X1536 N1536 N1537 Segment
X1537 N1537 N1538 Segment
X1538 N1538 N1539 Segment
X1539 N1539 N1540 Segment
X1540 N1540 N1541 Segment
X1541 N1541 N1542 Segment
X1542 N1542 N1543 Segment
X1543 N1543 N1544 Segment
X1544 N1544 N1545 Segment
X1545 N1545 N1546 Segment
X1546 N1546 N1547 Segment
X1547 N1547 N1548 Segment
X1548 N1548 N1549 Segment
X1549 N1549 N1550 Segment
X1550 N1550 N1551 Segment
X1551 N1551 N1552 Segment
X1552 N1552 N1553 Segment
X1553 N1553 N1554 Segment
X1554 N1554 N1555 Segment
X1555 N1555 N1556 Segment
X1556 N1556 N1557 Segment
X1557 N1557 N1558 Segment
X1558 N1558 N1559 Segment
X1559 N1559 N1560 Segment
X1560 N1560 N1561 Segment
X1561 N1561 N1562 Segment
X1562 N1562 N1563 Segment
X1563 N1563 N1564 Segment
X1564 N1564 N1565 Segment
X1565 N1565 N1566 Segment
X1566 N1566 N1567 Segment
X1567 N1567 N1568 Segment
X1568 N1568 N1569 Segment
X1569 N1569 N1570 Segment
X1570 N1570 N1571 Segment
X1571 N1571 N1572 Segment
X1572 N1572 N1573 Segment
X1573 N1573 N1574 Segment
X1574 N1574 N1575 Segment
X1575 N1575 N1576 Segment
X1576 N1576 N1577 Segment
X1577 N1577 N1578 Segment
X1578 N1578 N1579 Segment
X1579 N1579 N1580 Segment
X1580 N1580 N1581 Segment
X1581 N1581 N1582 Segment
X1582 N1582 N1583 Segment
X1583 N1583 N1584 Segment
X1584 N1584 N1585 Segment
X1585 N1585 N1586 Segment
X1586 N1586 N1587 Segment
X1587 N1587 N1588 Segment
X1588 N1588 N1589 Segment
X1589 N1589 N1590 Segment
X1590 N1590 N1591 Segment
X1591 N1591 N1592 Segment
X1592 N1592 N1593 Segment
X1593 N1593 N1594 Segment
X1594 N1594 N1595 Segment
X1595 N1595 N1596 Segment
X1596 N1596 N1597 Segment
X1597 N1597 N1598 Segment
X1598 N1598 N1599 Segment
X1599 N1599 N1600 Segment
X1600 N1600 N1601 Segment
X1601 N1601 N1602 Segment
X1602 N1602 N1603 Segment
X1603 N1603 N1604 Segment
X1604 N1604 N1605 Segment
X1605 N1605 N1606 Segment
X1606 N1606 N1607 Segment
X1607 N1607 N1608 Segment
X1608 N1608 N1609 Segment
X1609 N1609 N1610 Segment
X1610 N1610 N1611 Segment
X1611 N1611 N1612 Segment
X1612 N1612 N1613 Segment
X1613 N1613 N1614 Segment
X1614 N1614 N1615 Segment
X1615 N1615 N1616 Segment
X1616 N1616 N1617 Segment
X1617 N1617 N1618 Segment
X1618 N1618 N1619 Segment
X1619 N1619 N1620 Segment
X1620 N1620 N1621 Segment
X1621 N1621 N1622 Segment
X1622 N1622 N1623 Segment
X1623 N1623 N1624 Segment
X1624 N1624 N1625 Segment
X1625 N1625 N1626 Segment
X1626 N1626 N1627 Segment
X1627 N1627 N1628 Segment
X1628 N1628 N1629 Segment
X1629 N1629 N1630 Segment
X1630 N1630 N1631 Segment
X1631 N1631 N1632 Segment
X1632 N1632 N1633 Segment
X1633 N1633 N1634 Segment
X1634 N1634 N1635 Segment
X1635 N1635 N1636 Segment
X1636 N1636 N1637 Segment
X1637 N1637 N1638 Segment
X1638 N1638 N1639 Segment
X1639 N1639 N1640 Segment
X1640 N1640 N1641 Segment
X1641 N1641 N1642 Segment
X1642 N1642 N1643 Segment
X1643 N1643 N1644 Segment
X1644 N1644 N1645 Segment
X1645 N1645 N1646 Segment
X1646 N1646 N1647 Segment
X1647 N1647 N1648 Segment
X1648 N1648 N1649 Segment
X1649 N1649 N1650 Segment
X1650 N1650 N1651 Segment
X1651 N1651 N1652 Segment
X1652 N1652 N1653 Segment
X1653 N1653 N1654 Segment
X1654 N1654 N1655 Segment
X1655 N1655 N1656 Segment
X1656 N1656 N1657 Segment
X1657 N1657 N1658 Segment
X1658 N1658 N1659 Segment
X1659 N1659 N1660 Segment
X1660 N1660 N1661 Segment
X1661 N1661 N1662 Segment
X1662 N1662 N1663 Segment
X1663 N1663 N1664 Segment
X1664 N1664 N1665 Segment
X1665 N1665 N1666 Segment
X1666 N1666 N1667 Segment
X1667 N1667 N1668 Segment
X1668 N1668 N1669 Segment
X1669 N1669 N1670 Segment
X1670 N1670 N1671 Segment
X1671 N1671 N1672 Segment
X1672 N1672 N1673 Segment
X1673 N1673 N1674 Segment
X1674 N1674 N1675 Segment
X1675 N1675 N1676 Segment
X1676 N1676 N1677 Segment
X1677 N1677 N1678 Segment
X1678 N1678 N1679 Segment
X1679 N1679 N1680 Segment
X1680 N1680 N1681 Segment
X1681 N1681 N1682 Segment
X1682 N1682 N1683 Segment
X1683 N1683 N1684 Segment
X1684 N1684 N1685 Segment
X1685 N1685 N1686 Segment
X1686 N1686 N1687 Segment
X1687 N1687 N1688 Segment
X1688 N1688 N1689 Segment
X1689 N1689 N1690 Segment
X1690 N1690 N1691 Segment
X1691 N1691 N1692 Segment
X1692 N1692 N1693 Segment
X1693 N1693 N1694 Segment
X1694 N1694 N1695 Segment
X1695 N1695 N1696 Segment
X1696 N1696 N1697 Segment
X1697 N1697 N1698 Segment
X1698 N1698 N1699 Segment
X1699 N1699 N1700 Segment
X1700 N1700 N1701 Segment
X1701 N1701 N1702 Segment
X1702 N1702 N1703 Segment
X1703 N1703 N1704 Segment
X1704 N1704 N1705 Segment
X1705 N1705 N1706 Segment
X1706 N1706 N1707 Segment
X1707 N1707 N1708 Segment
X1708 N1708 N1709 Segment
X1709 N1709 N1710 Segment
X1710 N1710 N1711 Segment
X1711 N1711 N1712 Segment
X1712 N1712 N1713 Segment
X1713 N1713 N1714 Segment
X1714 N1714 N1715 Segment
X1715 N1715 N1716 Segment
X1716 N1716 N1717 Segment
X1717 N1717 N1718 Segment
X1718 N1718 N1719 Segment
X1719 N1719 N1720 Segment
X1720 N1720 N1721 Segment
X1721 N1721 N1722 Segment
X1722 N1722 N1723 Segment
X1723 N1723 N1724 Segment
X1724 N1724 N1725 Segment
X1725 N1725 N1726 Segment
X1726 N1726 N1727 Segment
X1727 N1727 N1728 Segment
X1728 N1728 N1729 Segment
X1729 N1729 N1730 Segment
X1730 N1730 N1731 Segment
X1731 N1731 N1732 Segment
X1732 N1732 N1733 Segment
X1733 N1733 N1734 Segment
X1734 N1734 N1735 Segment
X1735 N1735 N1736 Segment
X1736 N1736 N1737 Segment
X1737 N1737 N1738 Segment
X1738 N1738 N1739 Segment
X1739 N1739 N1740 Segment
X1740 N1740 N1741 Segment
X1741 N1741 N1742 Segment
X1742 N1742 N1743 Segment
X1743 N1743 N1744 Segment
X1744 N1744 N1745 Segment
X1745 N1745 N1746 Segment
X1746 N1746 N1747 Segment
X1747 N1747 N1748 Segment
X1748 N1748 N1749 Segment
X1749 N1749 N1750 Segment
X1750 N1750 N1751 Segment
X1751 N1751 N1752 Segment
X1752 N1752 N1753 Segment
X1753 N1753 N1754 Segment
X1754 N1754 N1755 Segment
X1755 N1755 N1756 Segment
X1756 N1756 N1757 Segment
X1757 N1757 N1758 Segment
X1758 N1758 N1759 Segment
X1759 N1759 N1760 Segment
X1760 N1760 N1761 Segment
X1761 N1761 N1762 Segment
X1762 N1762 N1763 Segment
X1763 N1763 N1764 Segment
X1764 N1764 N1765 Segment
X1765 N1765 N1766 Segment
X1766 N1766 N1767 Segment
X1767 N1767 N1768 Segment
X1768 N1768 N1769 Segment
X1769 N1769 N1770 Segment
X1770 N1770 N1771 Segment
X1771 N1771 N1772 Segment
X1772 N1772 N1773 Segment
X1773 N1773 N1774 Segment
X1774 N1774 N1775 Segment
X1775 N1775 N1776 Segment
X1776 N1776 N1777 Segment
X1777 N1777 N1778 Segment
X1778 N1778 N1779 Segment
X1779 N1779 N1780 Segment
X1780 N1780 N1781 Segment
X1781 N1781 N1782 Segment
X1782 N1782 N1783 Segment
X1783 N1783 N1784 Segment
X1784 N1784 N1785 Segment
X1785 N1785 N1786 Segment
X1786 N1786 N1787 Segment
X1787 N1787 N1788 Segment
X1788 N1788 N1789 Segment
X1789 N1789 N1790 Segment
X1790 N1790 N1791 Segment
X1791 N1791 N1792 Segment
X1792 N1792 N1793 Segment
X1793 N1793 N1794 Segment
X1794 N1794 N1795 Segment
X1795 N1795 N1796 Segment
X1796 N1796 N1797 Segment
X1797 N1797 N1798 Segment
X1798 N1798 N1799 Segment
X1799 N1799 N1800 Segment
X1800 N1800 N1801 Segment
X1801 N1801 N1802 Segment
X1802 N1802 N1803 Segment
X1803 N1803 N1804 Segment
X1804 N1804 N1805 Segment
X1805 N1805 N1806 Segment
X1806 N1806 N1807 Segment
X1807 N1807 N1808 Segment
X1808 N1808 N1809 Segment
X1809 N1809 N1810 Segment
X1810 N1810 N1811 Segment
X1811 N1811 N1812 Segment
X1812 N1812 N1813 Segment
X1813 N1813 N1814 Segment
X1814 N1814 N1815 Segment
X1815 N1815 N1816 Segment
X1816 N1816 N1817 Segment
X1817 N1817 N1818 Segment
X1818 N1818 N1819 Segment
X1819 N1819 N1820 Segment
X1820 N1820 N1821 Segment
X1821 N1821 N1822 Segment
X1822 N1822 N1823 Segment
X1823 N1823 N1824 Segment
X1824 N1824 N1825 Segment
X1825 N1825 N1826 Segment
X1826 N1826 N1827 Segment
X1827 N1827 N1828 Segment
X1828 N1828 N1829 Segment
X1829 N1829 N1830 Segment
X1830 N1830 N1831 Segment
X1831 N1831 N1832 Segment
X1832 N1832 N1833 Segment
X1833 N1833 N1834 Segment
X1834 N1834 N1835 Segment
X1835 N1835 N1836 Segment
X1836 N1836 N1837 Segment
X1837 N1837 N1838 Segment
X1838 N1838 N1839 Segment
X1839 N1839 N1840 Segment
X1840 N1840 N1841 Segment
X1841 N1841 N1842 Segment
X1842 N1842 N1843 Segment
X1843 N1843 N1844 Segment
X1844 N1844 N1845 Segment
X1845 N1845 N1846 Segment
X1846 N1846 N1847 Segment
X1847 N1847 N1848 Segment
X1848 N1848 N1849 Segment
X1849 N1849 N1850 Segment
X1850 N1850 N1851 Segment
X1851 N1851 N1852 Segment
X1852 N1852 N1853 Segment
X1853 N1853 N1854 Segment
X1854 N1854 N1855 Segment
X1855 N1855 N1856 Segment
X1856 N1856 N1857 Segment
X1857 N1857 N1858 Segment
X1858 N1858 N1859 Segment
X1859 N1859 N1860 Segment
X1860 N1860 N1861 Segment
X1861 N1861 N1862 Segment
X1862 N1862 N1863 Segment
X1863 N1863 N1864 Segment
X1864 N1864 N1865 Segment
X1865 N1865 N1866 Segment
X1866 N1866 N1867 Segment
X1867 N1867 N1868 Segment
X1868 N1868 N1869 Segment
X1869 N1869 N1870 Segment
X1870 N1870 N1871 Segment
X1871 N1871 N1872 Segment
X1872 N1872 N1873 Segment
X1873 N1873 N1874 Segment
X1874 N1874 N1875 Segment
X1875 N1875 N1876 Segment
X1876 N1876 N1877 Segment
X1877 N1877 N1878 Segment
X1878 N1878 N1879 Segment
X1879 N1879 N1880 Segment
X1880 N1880 N1881 Segment
X1881 N1881 N1882 Segment
X1882 N1882 N1883 Segment
X1883 N1883 N1884 Segment
X1884 N1884 N1885 Segment
X1885 N1885 N1886 Segment
X1886 N1886 N1887 Segment
X1887 N1887 N1888 Segment
X1888 N1888 N1889 Segment
X1889 N1889 N1890 Segment
X1890 N1890 N1891 Segment
X1891 N1891 N1892 Segment
X1892 N1892 N1893 Segment
X1893 N1893 N1894 Segment
X1894 N1894 N1895 Segment
X1895 N1895 N1896 Segment
X1896 N1896 N1897 Segment
X1897 N1897 N1898 Segment
X1898 N1898 N1899 Segment
X1899 N1899 N1900 Segment
X1900 N1900 N1901 Segment
X1901 N1901 N1902 Segment
X1902 N1902 N1903 Segment
X1903 N1903 N1904 Segment
X1904 N1904 N1905 Segment
X1905 N1905 N1906 Segment
X1906 N1906 N1907 Segment
X1907 N1907 N1908 Segment
X1908 N1908 N1909 Segment
X1909 N1909 N1910 Segment
X1910 N1910 N1911 Segment
X1911 N1911 N1912 Segment
X1912 N1912 N1913 Segment
X1913 N1913 N1914 Segment
X1914 N1914 N1915 Segment
X1915 N1915 N1916 Segment
X1916 N1916 N1917 Segment
X1917 N1917 N1918 Segment
X1918 N1918 N1919 Segment
X1919 N1919 N1920 Segment
X1920 N1920 N1921 Segment
X1921 N1921 N1922 Segment
X1922 N1922 N1923 Segment
X1923 N1923 N1924 Segment
X1924 N1924 N1925 Segment
X1925 N1925 N1926 Segment
X1926 N1926 N1927 Segment
X1927 N1927 N1928 Segment
X1928 N1928 N1929 Segment
X1929 N1929 N1930 Segment
X1930 N1930 N1931 Segment
X1931 N1931 N1932 Segment
X1932 N1932 N1933 Segment
X1933 N1933 N1934 Segment
X1934 N1934 N1935 Segment
X1935 N1935 N1936 Segment
X1936 N1936 N1937 Segment
X1937 N1937 N1938 Segment
X1938 N1938 N1939 Segment
X1939 N1939 N1940 Segment
X1940 N1940 N1941 Segment
X1941 N1941 N1942 Segment
X1942 N1942 N1943 Segment
X1943 N1943 N1944 Segment
X1944 N1944 N1945 Segment
X1945 N1945 N1946 Segment
X1946 N1946 N1947 Segment
X1947 N1947 N1948 Segment
X1948 N1948 N1949 Segment
X1949 N1949 N1950 Segment
X1950 N1950 N1951 Segment
X1951 N1951 N1952 Segment
X1952 N1952 N1953 Segment
X1953 N1953 N1954 Segment
X1954 N1954 N1955 Segment
X1955 N1955 N1956 Segment
X1956 N1956 N1957 Segment
X1957 N1957 N1958 Segment
X1958 N1958 N1959 Segment
X1959 N1959 N1960 Segment
X1960 N1960 N1961 Segment
X1961 N1961 N1962 Segment
X1962 N1962 N1963 Segment
X1963 N1963 N1964 Segment
X1964 N1964 N1965 Segment
X1965 N1965 N1966 Segment
X1966 N1966 N1967 Segment
X1967 N1967 N1968 Segment
X1968 N1968 N1969 Segment
X1969 N1969 N1970 Segment
X1970 N1970 N1971 Segment
X1971 N1971 N1972 Segment
X1972 N1972 N1973 Segment
X1973 N1973 N1974 Segment
X1974 N1974 N1975 Segment
X1975 N1975 N1976 Segment
X1976 N1976 N1977 Segment
X1977 N1977 N1978 Segment
X1978 N1978 N1979 Segment
X1979 N1979 N1980 Segment
X1980 N1980 N1981 Segment
X1981 N1981 N1982 Segment
X1982 N1982 N1983 Segment
X1983 N1983 N1984 Segment
X1984 N1984 N1985 Segment
X1985 N1985 N1986 Segment
X1986 N1986 N1987 Segment
X1987 N1987 N1988 Segment
X1988 N1988 N1989 Segment
X1989 N1989 N1990 Segment
X1990 N1990 N1991 Segment
X1991 N1991 N1992 Segment
X1992 N1992 N1993 Segment
X1993 N1993 N1994 Segment
X1994 N1994 N1995 Segment
X1995 N1995 N1996 Segment
X1996 N1996 N1997 Segment
X1997 N1997 N1998 Segment
X1998 N1998 N1999 Segment
X1999 N1999 N2000 Segment
X2000 N2000 N2001 Segment
X2001 N2001 N2002 Segment
X2002 N2002 N2003 Segment
X2003 N2003 N2004 Segment
X2004 N2004 N2005 Segment
X2005 N2005 N2006 Segment
X2006 N2006 N2007 Segment
X2007 N2007 N2008 Segment
X2008 N2008 N2009 Segment
X2009 N2009 N2010 Segment
X2010 N2010 N2011 Segment
X2011 N2011 N2012 Segment
X2012 N2012 N2013 Segment
X2013 N2013 N2014 Segment
X2014 N2014 N2015 Segment
X2015 N2015 N2016 Segment
X2016 N2016 N2017 Segment
X2017 N2017 N2018 Segment
X2018 N2018 N2019 Segment
X2019 N2019 N2020 Segment
X2020 N2020 N2021 Segment
X2021 N2021 N2022 Segment
X2022 N2022 N2023 Segment
X2023 N2023 N2024 Segment
X2024 N2024 N2025 Segment
X2025 N2025 N2026 Segment
X2026 N2026 N2027 Segment
X2027 N2027 N2028 Segment
X2028 N2028 N2029 Segment
X2029 N2029 N2030 Segment
X2030 N2030 N2031 Segment
X2031 N2031 N2032 Segment
X2032 N2032 N2033 Segment
X2033 N2033 N2034 Segment
X2034 N2034 N2035 Segment
X2035 N2035 N2036 Segment
X2036 N2036 N2037 Segment
X2037 N2037 N2038 Segment
X2038 N2038 N2039 Segment
X2039 N2039 N2040 Segment
X2040 N2040 N2041 Segment
X2041 N2041 N2042 Segment
X2042 N2042 N2043 Segment
X2043 N2043 N2044 Segment
X2044 N2044 N2045 Segment
X2045 N2045 N2046 Segment
X2046 N2046 N2047 Segment
X2047 N2047 N2048 Segment
X2048 N2048 N2049 Segment
X2049 N2049 N2050 Segment
X2050 N2050 N2051 Segment
X2051 N2051 N2052 Segment
X2052 N2052 N2053 Segment
X2053 N2053 N2054 Segment
X2054 N2054 N2055 Segment
X2055 N2055 N2056 Segment
X2056 N2056 N2057 Segment
X2057 N2057 N2058 Segment
X2058 N2058 N2059 Segment
X2059 N2059 N2060 Segment
X2060 N2060 N2061 Segment
X2061 N2061 N2062 Segment
X2062 N2062 N2063 Segment
X2063 N2063 N2064 Segment
X2064 N2064 N2065 Segment
X2065 N2065 N2066 Segment
X2066 N2066 N2067 Segment
X2067 N2067 N2068 Segment
X2068 N2068 N2069 Segment
X2069 N2069 N2070 Segment
X2070 N2070 N2071 Segment
X2071 N2071 N2072 Segment
X2072 N2072 N2073 Segment
X2073 N2073 N2074 Segment
X2074 N2074 N2075 Segment
X2075 N2075 N2076 Segment
X2076 N2076 N2077 Segment
X2077 N2077 N2078 Segment
X2078 N2078 N2079 Segment
X2079 N2079 N2080 Segment
X2080 N2080 N2081 Segment
X2081 N2081 N2082 Segment
X2082 N2082 N2083 Segment
X2083 N2083 N2084 Segment
X2084 N2084 N2085 Segment
X2085 N2085 N2086 Segment
X2086 N2086 N2087 Segment
X2087 N2087 N2088 Segment
X2088 N2088 N2089 Segment
X2089 N2089 N2090 Segment
X2090 N2090 N2091 Segment
X2091 N2091 N2092 Segment
X2092 N2092 N2093 Segment
X2093 N2093 N2094 Segment
X2094 N2094 N2095 Segment
X2095 N2095 N2096 Segment
X2096 N2096 N2097 Segment
X2097 N2097 N2098 Segment
X2098 N2098 N2099 Segment
X2099 N2099 N2100 Segment
X2100 N2100 N2101 Segment
X2101 N2101 N2102 Segment
X2102 N2102 N2103 Segment
X2103 N2103 N2104 Segment
X2104 N2104 N2105 Segment
X2105 N2105 N2106 Segment
X2106 N2106 N2107 Segment
X2107 N2107 N2108 Segment
X2108 N2108 N2109 Segment
X2109 N2109 N2110 Segment
X2110 N2110 N2111 Segment
X2111 N2111 N2112 Segment
X2112 N2112 N2113 Segment
X2113 N2113 N2114 Segment
X2114 N2114 N2115 Segment
X2115 N2115 N2116 Segment
X2116 N2116 N2117 Segment
X2117 N2117 N2118 Segment
X2118 N2118 N2119 Segment
X2119 N2119 N2120 Segment
X2120 N2120 N2121 Segment
X2121 N2121 N2122 Segment
X2122 N2122 N2123 Segment
X2123 N2123 N2124 Segment
X2124 N2124 N2125 Segment
X2125 N2125 N2126 Segment
X2126 N2126 N2127 Segment
X2127 N2127 N2128 Segment
X2128 N2128 N2129 Segment
X2129 N2129 N2130 Segment
X2130 N2130 N2131 Segment
X2131 N2131 N2132 Segment
X2132 N2132 N2133 Segment
X2133 N2133 N2134 Segment
X2134 N2134 N2135 Segment
X2135 N2135 N2136 Segment
X2136 N2136 N2137 Segment
X2137 N2137 N2138 Segment
X2138 N2138 N2139 Segment
X2139 N2139 N2140 Segment
X2140 N2140 N2141 Segment
X2141 N2141 N2142 Segment
X2142 N2142 N2143 Segment
X2143 N2143 N2144 Segment
X2144 N2144 N2145 Segment
X2145 N2145 N2146 Segment
X2146 N2146 N2147 Segment
X2147 N2147 N2148 Segment
X2148 N2148 N2149 Segment
X2149 N2149 N2150 Segment
X2150 N2150 N2151 Segment
X2151 N2151 N2152 Segment
X2152 N2152 N2153 Segment
X2153 N2153 N2154 Segment
X2154 N2154 N2155 Segment
X2155 N2155 N2156 Segment
X2156 N2156 N2157 Segment
X2157 N2157 N2158 Segment
X2158 N2158 N2159 Segment
X2159 N2159 N2160 Segment
X2160 N2160 N2161 Segment
X2161 N2161 N2162 Segment
X2162 N2162 N2163 Segment
X2163 N2163 N2164 Segment
X2164 N2164 N2165 Segment
X2165 N2165 N2166 Segment
X2166 N2166 N2167 Segment
X2167 N2167 N2168 Segment
X2168 N2168 N2169 Segment
X2169 N2169 N2170 Segment
X2170 N2170 N2171 Segment
X2171 N2171 N2172 Segment
X2172 N2172 N2173 Segment
X2173 N2173 N2174 Segment
X2174 N2174 N2175 Segment
X2175 N2175 N2176 Segment
X2176 N2176 N2177 Segment
X2177 N2177 N2178 Segment
X2178 N2178 N2179 Segment
X2179 N2179 N2180 Segment
X2180 N2180 N2181 Segment
X2181 N2181 N2182 Segment
X2182 N2182 N2183 Segment
X2183 N2183 N2184 Segment
X2184 N2184 N2185 Segment
X2185 N2185 N2186 Segment
X2186 N2186 N2187 Segment
X2187 N2187 N2188 Segment
X2188 N2188 N2189 Segment
X2189 N2189 N2190 Segment
X2190 N2190 N2191 Segment
X2191 N2191 N2192 Segment
X2192 N2192 N2193 Segment
X2193 N2193 N2194 Segment
X2194 N2194 N2195 Segment
X2195 N2195 N2196 Segment
X2196 N2196 N2197 Segment
X2197 N2197 N2198 Segment
X2198 N2198 N2199 Segment
X2199 N2199 N2200 Segment
X2200 N2200 N2201 Segment
X2201 N2201 N2202 Segment
X2202 N2202 N2203 Segment
X2203 N2203 N2204 Segment
X2204 N2204 N2205 Segment
X2205 N2205 N2206 Segment
X2206 N2206 N2207 Segment
X2207 N2207 N2208 Segment
X2208 N2208 N2209 Segment
X2209 N2209 N2210 Segment
X2210 N2210 N2211 Segment
X2211 N2211 N2212 Segment
X2212 N2212 N2213 Segment
X2213 N2213 N2214 Segment
X2214 N2214 N2215 Segment
X2215 N2215 N2216 Segment
X2216 N2216 N2217 Segment
X2217 N2217 N2218 Segment
X2218 N2218 N2219 Segment
X2219 N2219 N2220 Segment
X2220 N2220 N2221 Segment
X2221 N2221 N2222 Segment
X2222 N2222 N2223 Segment
X2223 N2223 N2224 Segment
X2224 N2224 N2225 Segment
X2225 N2225 N2226 Segment
X2226 N2226 N2227 Segment
X2227 N2227 N2228 Segment
X2228 N2228 N2229 Segment
X2229 N2229 N2230 Segment
X2230 N2230 N2231 Segment
X2231 N2231 N2232 Segment
X2232 N2232 N2233 Segment
X2233 N2233 N2234 Segment
X2234 N2234 N2235 Segment
X2235 N2235 N2236 Segment
X2236 N2236 N2237 Segment
X2237 N2237 N2238 Segment
X2238 N2238 N2239 Segment
X2239 N2239 N2240 Segment
X2240 N2240 N2241 Segment
X2241 N2241 N2242 Segment
X2242 N2242 N2243 Segment
X2243 N2243 N2244 Segment
X2244 N2244 N2245 Segment
X2245 N2245 N2246 Segment
X2246 N2246 N2247 Segment
X2247 N2247 N2248 Segment
X2248 N2248 N2249 Segment
X2249 N2249 N2250 Segment
X2250 N2250 N2251 Segment
X2251 N2251 N2252 Segment
X2252 N2252 N2253 Segment
X2253 N2253 N2254 Segment
X2254 N2254 N2255 Segment
X2255 N2255 N2256 Segment
X2256 N2256 N2257 Segment
X2257 N2257 N2258 Segment
X2258 N2258 N2259 Segment
X2259 N2259 N2260 Segment
X2260 N2260 N2261 Segment
X2261 N2261 N2262 Segment
X2262 N2262 N2263 Segment
X2263 N2263 N2264 Segment
X2264 N2264 N2265 Segment
X2265 N2265 N2266 Segment
X2266 N2266 N2267 Segment
X2267 N2267 N2268 Segment
X2268 N2268 N2269 Segment
X2269 N2269 N2270 Segment
X2270 N2270 N2271 Segment
X2271 N2271 N2272 Segment
X2272 N2272 N2273 Segment
X2273 N2273 N2274 Segment
X2274 N2274 N2275 Segment
X2275 N2275 N2276 Segment
X2276 N2276 N2277 Segment
X2277 N2277 N2278 Segment
X2278 N2278 N2279 Segment
X2279 N2279 N2280 Segment
X2280 N2280 N2281 Segment
X2281 N2281 N2282 Segment
X2282 N2282 N2283 Segment
X2283 N2283 N2284 Segment
X2284 N2284 N2285 Segment
X2285 N2285 N2286 Segment
X2286 N2286 N2287 Segment
X2287 N2287 N2288 Segment
X2288 N2288 N2289 Segment
X2289 N2289 N2290 Segment
X2290 N2290 N2291 Segment
X2291 N2291 N2292 Segment
X2292 N2292 N2293 Segment
X2293 N2293 N2294 Segment
X2294 N2294 N2295 Segment
X2295 N2295 N2296 Segment
X2296 N2296 N2297 Segment
X2297 N2297 N2298 Segment
X2298 N2298 N2299 Segment
X2299 N2299 N2300 Segment
X2300 N2300 N2301 Segment
X2301 N2301 N2302 Segment
X2302 N2302 N2303 Segment
X2303 N2303 N2304 Segment
X2304 N2304 N2305 Segment
X2305 N2305 N2306 Segment
X2306 N2306 N2307 Segment
X2307 N2307 N2308 Segment
X2308 N2308 N2309 Segment
X2309 N2309 N2310 Segment
X2310 N2310 N2311 Segment
X2311 N2311 N2312 Segment
X2312 N2312 N2313 Segment
X2313 N2313 N2314 Segment
X2314 N2314 N2315 Segment
X2315 N2315 N2316 Segment
X2316 N2316 N2317 Segment
X2317 N2317 N2318 Segment
X2318 N2318 N2319 Segment
X2319 N2319 N2320 Segment
X2320 N2320 N2321 Segment
X2321 N2321 N2322 Segment
X2322 N2322 N2323 Segment
X2323 N2323 N2324 Segment
X2324 N2324 N2325 Segment
X2325 N2325 N2326 Segment
X2326 N2326 N2327 Segment
X2327 N2327 N2328 Segment
X2328 N2328 N2329 Segment
X2329 N2329 N2330 Segment
X2330 N2330 N2331 Segment
X2331 N2331 N2332 Segment
X2332 N2332 N2333 Segment
X2333 N2333 N2334 Segment
X2334 N2334 N2335 Segment
X2335 N2335 N2336 Segment
X2336 N2336 N2337 Segment
X2337 N2337 N2338 Segment
X2338 N2338 N2339 Segment
X2339 N2339 N2340 Segment
X2340 N2340 N2341 Segment
X2341 N2341 N2342 Segment
X2342 N2342 N2343 Segment
X2343 N2343 N2344 Segment
X2344 N2344 N2345 Segment
X2345 N2345 N2346 Segment
X2346 N2346 N2347 Segment
X2347 N2347 N2348 Segment
X2348 N2348 N2349 Segment
X2349 N2349 N2350 Segment
X2350 N2350 N2351 Segment
X2351 N2351 N2352 Segment
X2352 N2352 N2353 Segment
X2353 N2353 N2354 Segment
X2354 N2354 N2355 Segment
X2355 N2355 N2356 Segment
X2356 N2356 N2357 Segment
X2357 N2357 N2358 Segment
X2358 N2358 N2359 Segment
X2359 N2359 N2360 Segment
X2360 N2360 N2361 Segment
X2361 N2361 N2362 Segment
X2362 N2362 N2363 Segment
X2363 N2363 N2364 Segment
X2364 N2364 N2365 Segment
X2365 N2365 N2366 Segment
X2366 N2366 N2367 Segment
X2367 N2367 N2368 Segment
X2368 N2368 N2369 Segment
X2369 N2369 N2370 Segment
X2370 N2370 N2371 Segment
X2371 N2371 N2372 Segment
X2372 N2372 N2373 Segment
X2373 N2373 N2374 Segment
X2374 N2374 N2375 Segment
X2375 N2375 N2376 Segment
X2376 N2376 N2377 Segment
X2377 N2377 N2378 Segment
X2378 N2378 N2379 Segment
X2379 N2379 N2380 Segment
X2380 N2380 N2381 Segment
X2381 N2381 N2382 Segment
X2382 N2382 N2383 Segment
X2383 N2383 N2384 Segment
X2384 N2384 N2385 Segment
X2385 N2385 N2386 Segment
X2386 N2386 N2387 Segment
X2387 N2387 N2388 Segment
X2388 N2388 N2389 Segment
X2389 N2389 N2390 Segment
X2390 N2390 N2391 Segment
X2391 N2391 N2392 Segment
X2392 N2392 N2393 Segment
X2393 N2393 N2394 Segment
X2394 N2394 N2395 Segment
X2395 N2395 N2396 Segment
X2396 N2396 N2397 Segment
X2397 N2397 N2398 Segment
X2398 N2398 N2399 Segment
X2399 N2399 N2400 Segment
X2400 N2400 N2401 Segment
X2401 N2401 N2402 Segment
X2402 N2402 N2403 Segment
X2403 N2403 N2404 Segment
X2404 N2404 N2405 Segment
X2405 N2405 N2406 Segment
X2406 N2406 N2407 Segment
X2407 N2407 N2408 Segment
X2408 N2408 N2409 Segment
X2409 N2409 N2410 Segment
X2410 N2410 N2411 Segment
X2411 N2411 N2412 Segment
X2412 N2412 N2413 Segment
X2413 N2413 N2414 Segment
X2414 N2414 N2415 Segment
X2415 N2415 N2416 Segment
X2416 N2416 N2417 Segment
X2417 N2417 N2418 Segment
X2418 N2418 N2419 Segment
X2419 N2419 N2420 Segment
X2420 N2420 N2421 Segment
X2421 N2421 N2422 Segment
X2422 N2422 N2423 Segment
X2423 N2423 N2424 Segment
X2424 N2424 N2425 Segment
X2425 N2425 N2426 Segment
X2426 N2426 N2427 Segment
X2427 N2427 N2428 Segment
X2428 N2428 N2429 Segment
X2429 N2429 N2430 Segment
X2430 N2430 N2431 Segment
X2431 N2431 N2432 Segment
X2432 N2432 N2433 Segment
X2433 N2433 N2434 Segment
X2434 N2434 N2435 Segment
X2435 N2435 N2436 Segment
X2436 N2436 N2437 Segment
X2437 N2437 N2438 Segment
X2438 N2438 N2439 Segment
X2439 N2439 N2440 Segment
X2440 N2440 N2441 Segment
X2441 N2441 N2442 Segment
X2442 N2442 N2443 Segment
X2443 N2443 N2444 Segment
X2444 N2444 N2445 Segment
X2445 N2445 N2446 Segment
X2446 N2446 N2447 Segment
X2447 N2447 N2448 Segment
X2448 N2448 N2449 Segment
X2449 N2449 N2450 Segment
X2450 N2450 N2451 Segment
X2451 N2451 N2452 Segment
X2452 N2452 N2453 Segment
X2453 N2453 N2454 Segment
X2454 N2454 N2455 Segment
X2455 N2455 N2456 Segment
X2456 N2456 N2457 Segment
X2457 N2457 N2458 Segment
X2458 N2458 N2459 Segment
X2459 N2459 N2460 Segment
X2460 N2460 N2461 Segment
X2461 N2461 N2462 Segment
X2462 N2462 N2463 Segment
X2463 N2463 N2464 Segment
X2464 N2464 N2465 Segment
X2465 N2465 N2466 Segment
X2466 N2466 N2467 Segment
X2467 N2467 N2468 Segment
X2468 N2468 N2469 Segment
X2469 N2469 N2470 Segment
X2470 N2470 N2471 Segment
X2471 N2471 N2472 Segment
X2472 N2472 N2473 Segment
X2473 N2473 N2474 Segment
X2474 N2474 N2475 Segment
X2475 N2475 N2476 Segment
X2476 N2476 N2477 Segment
X2477 N2477 N2478 Segment
X2478 N2478 N2479 Segment
X2479 N2479 N2480 Segment
X2480 N2480 N2481 Segment
X2481 N2481 N2482 Segment
X2482 N2482 N2483 Segment
X2483 N2483 N2484 Segment
X2484 N2484 N2485 Segment
X2485 N2485 N2486 Segment
X2486 N2486 N2487 Segment
X2487 N2487 N2488 Segment
X2488 N2488 N2489 Segment
X2489 N2489 N2490 Segment
X2490 N2490 N2491 Segment
X2491 N2491 N2492 Segment
X2492 N2492 N2493 Segment
X2493 N2493 N2494 Segment
X2494 N2494 N2495 Segment
X2495 N2495 N2496 Segment
X2496 N2496 N2497 Segment
X2497 N2497 N2498 Segment
X2498 N2498 N2499 Segment
X2499 N2499 N2500 Segment
X2500 N2500 N2501 Segment
X2501 N2501 N2502 Segment
X2502 N2502 N2503 Segment
X2503 N2503 N2504 Segment
X2504 N2504 N2505 Segment
X2505 N2505 N2506 Segment
X2506 N2506 N2507 Segment
X2507 N2507 N2508 Segment
X2508 N2508 N2509 Segment
X2509 N2509 N2510 Segment
X2510 N2510 N2511 Segment
X2511 N2511 N2512 Segment
X2512 N2512 N2513 Segment
X2513 N2513 N2514 Segment
X2514 N2514 N2515 Segment
X2515 N2515 N2516 Segment
X2516 N2516 N2517 Segment
X2517 N2517 N2518 Segment
X2518 N2518 N2519 Segment
X2519 N2519 N2520 Segment
X2520 N2520 N2521 Segment
X2521 N2521 N2522 Segment
X2522 N2522 N2523 Segment
X2523 N2523 N2524 Segment
X2524 N2524 N2525 Segment
X2525 N2525 N2526 Segment
X2526 N2526 N2527 Segment
X2527 N2527 N2528 Segment
X2528 N2528 N2529 Segment
X2529 N2529 N2530 Segment
X2530 N2530 N2531 Segment
X2531 N2531 N2532 Segment
X2532 N2532 N2533 Segment
X2533 N2533 N2534 Segment
X2534 N2534 N2535 Segment
X2535 N2535 N2536 Segment
X2536 N2536 N2537 Segment
X2537 N2537 N2538 Segment
X2538 N2538 N2539 Segment
X2539 N2539 N2540 Segment
X2540 N2540 N2541 Segment
X2541 N2541 N2542 Segment
X2542 N2542 N2543 Segment
X2543 N2543 N2544 Segment
X2544 N2544 N2545 Segment
X2545 N2545 N2546 Segment
X2546 N2546 N2547 Segment
X2547 N2547 N2548 Segment
X2548 N2548 N2549 Segment
X2549 N2549 N2550 Segment
X2550 N2550 N2551 Segment
X2551 N2551 N2552 Segment
X2552 N2552 N2553 Segment
X2553 N2553 N2554 Segment
X2554 N2554 N2555 Segment
X2555 N2555 N2556 Segment
X2556 N2556 N2557 Segment
X2557 N2557 N2558 Segment
X2558 N2558 N2559 Segment
X2559 N2559 N2560 Segment
X2560 N2560 N2561 Segment
X2561 N2561 N2562 Segment
X2562 N2562 N2563 Segment
X2563 N2563 N2564 Segment
X2564 N2564 N2565 Segment
X2565 N2565 N2566 Segment
X2566 N2566 N2567 Segment
X2567 N2567 N2568 Segment
X2568 N2568 N2569 Segment
X2569 N2569 N2570 Segment
X2570 N2570 N2571 Segment
X2571 N2571 N2572 Segment
X2572 N2572 N2573 Segment
X2573 N2573 N2574 Segment
X2574 N2574 N2575 Segment
X2575 N2575 N2576 Segment
X2576 N2576 N2577 Segment
X2577 N2577 N2578 Segment
X2578 N2578 N2579 Segment
X2579 N2579 N2580 Segment
X2580 N2580 N2581 Segment
X2581 N2581 N2582 Segment
X2582 N2582 N2583 Segment
X2583 N2583 N2584 Segment
X2584 N2584 N2585 Segment
X2585 N2585 N2586 Segment
X2586 N2586 N2587 Segment
X2587 N2587 N2588 Segment
X2588 N2588 N2589 Segment
X2589 N2589 N2590 Segment
X2590 N2590 N2591 Segment
X2591 N2591 N2592 Segment
X2592 N2592 N2593 Segment
X2593 N2593 N2594 Segment
X2594 N2594 N2595 Segment
X2595 N2595 N2596 Segment
X2596 N2596 N2597 Segment
X2597 N2597 N2598 Segment
X2598 N2598 N2599 Segment
X2599 N2599 N2600 Segment
X2600 N2600 N2601 Segment
X2601 N2601 N2602 Segment
X2602 N2602 N2603 Segment
X2603 N2603 N2604 Segment
X2604 N2604 N2605 Segment
X2605 N2605 N2606 Segment
X2606 N2606 N2607 Segment
X2607 N2607 N2608 Segment
X2608 N2608 N2609 Segment
X2609 N2609 N2610 Segment
X2610 N2610 N2611 Segment
X2611 N2611 N2612 Segment
X2612 N2612 N2613 Segment
X2613 N2613 N2614 Segment
X2614 N2614 N2615 Segment
X2615 N2615 N2616 Segment
X2616 N2616 N2617 Segment
X2617 N2617 N2618 Segment
X2618 N2618 N2619 Segment
X2619 N2619 N2620 Segment
X2620 N2620 N2621 Segment
X2621 N2621 N2622 Segment
X2622 N2622 N2623 Segment
X2623 N2623 N2624 Segment
X2624 N2624 N2625 Segment
X2625 N2625 N2626 Segment
X2626 N2626 N2627 Segment
X2627 N2627 N2628 Segment
X2628 N2628 N2629 Segment
X2629 N2629 N2630 Segment
X2630 N2630 N2631 Segment
X2631 N2631 N2632 Segment
X2632 N2632 N2633 Segment
X2633 N2633 N2634 Segment
X2634 N2634 N2635 Segment
X2635 N2635 N2636 Segment
X2636 N2636 N2637 Segment
X2637 N2637 N2638 Segment
X2638 N2638 N2639 Segment
X2639 N2639 N2640 Segment
X2640 N2640 N2641 Segment
X2641 N2641 N2642 Segment
X2642 N2642 N2643 Segment
X2643 N2643 N2644 Segment
X2644 N2644 N2645 Segment
X2645 N2645 N2646 Segment
X2646 N2646 N2647 Segment
X2647 N2647 N2648 Segment
X2648 N2648 N2649 Segment
X2649 N2649 N2650 Segment
X2650 N2650 N2651 Segment
X2651 N2651 N2652 Segment
X2652 N2652 N2653 Segment
X2653 N2653 N2654 Segment
X2654 N2654 N2655 Segment
X2655 N2655 N2656 Segment
X2656 N2656 N2657 Segment
X2657 N2657 N2658 Segment
X2658 N2658 N2659 Segment
X2659 N2659 N2660 Segment
X2660 N2660 N2661 Segment
X2661 N2661 N2662 Segment
X2662 N2662 N2663 Segment
X2663 N2663 N2664 Segment
X2664 N2664 N2665 Segment
X2665 N2665 N2666 Segment
X2666 N2666 N2667 Segment
X2667 N2667 N2668 Segment
X2668 N2668 N2669 Segment
X2669 N2669 N2670 Segment
X2670 N2670 N2671 Segment
X2671 N2671 N2672 Segment
X2672 N2672 N2673 Segment
X2673 N2673 N2674 Segment
X2674 N2674 N2675 Segment
X2675 N2675 N2676 Segment
X2676 N2676 N2677 Segment
X2677 N2677 N2678 Segment
X2678 N2678 N2679 Segment
X2679 N2679 N2680 Segment
X2680 N2680 N2681 Segment
X2681 N2681 N2682 Segment
X2682 N2682 N2683 Segment
X2683 N2683 N2684 Segment
X2684 N2684 N2685 Segment
X2685 N2685 N2686 Segment
X2686 N2686 N2687 Segment
X2687 N2687 N2688 Segment
X2688 N2688 N2689 Segment
X2689 N2689 N2690 Segment
X2690 N2690 N2691 Segment
X2691 N2691 N2692 Segment
X2692 N2692 N2693 Segment
X2693 N2693 N2694 Segment
X2694 N2694 N2695 Segment
X2695 N2695 N2696 Segment
X2696 N2696 N2697 Segment
X2697 N2697 N2698 Segment
X2698 N2698 N2699 Segment
X2699 N2699 N2700 Segment
X2700 N2700 N2701 Segment
X2701 N2701 N2702 Segment
X2702 N2702 N2703 Segment
X2703 N2703 N2704 Segment
X2704 N2704 N2705 Segment
X2705 N2705 N2706 Segment
X2706 N2706 N2707 Segment
X2707 N2707 N2708 Segment
X2708 N2708 N2709 Segment
X2709 N2709 N2710 Segment
X2710 N2710 N2711 Segment
X2711 N2711 N2712 Segment
X2712 N2712 N2713 Segment
X2713 N2713 N2714 Segment
X2714 N2714 N2715 Segment
X2715 N2715 N2716 Segment
X2716 N2716 N2717 Segment
X2717 N2717 N2718 Segment
X2718 N2718 N2719 Segment
X2719 N2719 N2720 Segment
X2720 N2720 N2721 Segment
X2721 N2721 N2722 Segment
X2722 N2722 N2723 Segment
X2723 N2723 N2724 Segment
X2724 N2724 N2725 Segment
X2725 N2725 N2726 Segment
X2726 N2726 N2727 Segment
X2727 N2727 N2728 Segment
X2728 N2728 N2729 Segment
X2729 N2729 N2730 Segment
X2730 N2730 N2731 Segment
X2731 N2731 N2732 Segment
X2732 N2732 N2733 Segment
X2733 N2733 N2734 Segment
X2734 N2734 N2735 Segment
X2735 N2735 N2736 Segment
X2736 N2736 N2737 Segment
X2737 N2737 N2738 Segment
X2738 N2738 N2739 Segment
X2739 N2739 N2740 Segment
X2740 N2740 N2741 Segment
X2741 N2741 N2742 Segment
X2742 N2742 N2743 Segment
X2743 N2743 N2744 Segment
X2744 N2744 N2745 Segment
X2745 N2745 N2746 Segment
X2746 N2746 N2747 Segment
X2747 N2747 N2748 Segment
X2748 N2748 N2749 Segment
X2749 N2749 N2750 Segment
X2750 N2750 N2751 Segment
X2751 N2751 N2752 Segment
X2752 N2752 N2753 Segment
X2753 N2753 N2754 Segment
X2754 N2754 N2755 Segment
X2755 N2755 N2756 Segment
X2756 N2756 N2757 Segment
X2757 N2757 N2758 Segment
X2758 N2758 N2759 Segment
X2759 N2759 N2760 Segment
X2760 N2760 N2761 Segment
X2761 N2761 N2762 Segment
X2762 N2762 N2763 Segment
X2763 N2763 N2764 Segment
X2764 N2764 N2765 Segment
X2765 N2765 N2766 Segment
X2766 N2766 N2767 Segment
X2767 N2767 N2768 Segment
X2768 N2768 N2769 Segment
X2769 N2769 N2770 Segment
X2770 N2770 N2771 Segment
X2771 N2771 N2772 Segment
X2772 N2772 N2773 Segment
X2773 N2773 N2774 Segment
X2774 N2774 N2775 Segment
X2775 N2775 N2776 Segment
X2776 N2776 N2777 Segment
X2777 N2777 N2778 Segment
X2778 N2778 N2779 Segment
X2779 N2779 N2780 Segment
X2780 N2780 N2781 Segment
X2781 N2781 N2782 Segment
X2782 N2782 N2783 Segment
X2783 N2783 N2784 Segment
X2784 N2784 N2785 Segment
X2785 N2785 N2786 Segment
X2786 N2786 N2787 Segment
X2787 N2787 N2788 Segment
X2788 N2788 N2789 Segment
X2789 N2789 N2790 Segment
X2790 N2790 N2791 Segment
X2791 N2791 N2792 Segment
X2792 N2792 N2793 Segment
X2793 N2793 N2794 Segment
X2794 N2794 N2795 Segment
X2795 N2795 N2796 Segment
X2796 N2796 N2797 Segment
X2797 N2797 N2798 Segment
X2798 N2798 N2799 Segment
X2799 N2799 N2800 Segment
X2800 N2800 N2801 Segment
X2801 N2801 N2802 Segment
X2802 N2802 N2803 Segment
X2803 N2803 N2804 Segment
X2804 N2804 N2805 Segment
X2805 N2805 N2806 Segment
X2806 N2806 N2807 Segment
X2807 N2807 N2808 Segment
X2808 N2808 N2809 Segment
X2809 N2809 N2810 Segment
X2810 N2810 N2811 Segment
X2811 N2811 N2812 Segment
X2812 N2812 N2813 Segment
X2813 N2813 N2814 Segment
X2814 N2814 N2815 Segment
X2815 N2815 N2816 Segment
X2816 N2816 N2817 Segment
X2817 N2817 N2818 Segment
X2818 N2818 N2819 Segment
X2819 N2819 N2820 Segment
X2820 N2820 N2821 Segment
X2821 N2821 N2822 Segment
X2822 N2822 N2823 Segment
X2823 N2823 N2824 Segment
X2824 N2824 N2825 Segment
X2825 N2825 N2826 Segment
X2826 N2826 N2827 Segment
X2827 N2827 N2828 Segment
X2828 N2828 N2829 Segment
X2829 N2829 N2830 Segment
X2830 N2830 N2831 Segment
X2831 N2831 N2832 Segment
X2832 N2832 N2833 Segment
X2833 N2833 N2834 Segment
X2834 N2834 N2835 Segment
X2835 N2835 N2836 Segment
X2836 N2836 N2837 Segment
X2837 N2837 N2838 Segment
X2838 N2838 N2839 Segment
X2839 N2839 N2840 Segment
X2840 N2840 N2841 Segment
X2841 N2841 N2842 Segment
X2842 N2842 N2843 Segment
X2843 N2843 N2844 Segment
X2844 N2844 N2845 Segment
X2845 N2845 N2846 Segment
X2846 N2846 N2847 Segment
X2847 N2847 N2848 Segment
X2848 N2848 N2849 Segment
X2849 N2849 N2850 Segment
X2850 N2850 N2851 Segment
X2851 N2851 N2852 Segment
X2852 N2852 N2853 Segment
X2853 N2853 N2854 Segment
X2854 N2854 N2855 Segment
X2855 N2855 N2856 Segment
X2856 N2856 N2857 Segment
X2857 N2857 N2858 Segment
X2858 N2858 N2859 Segment
X2859 N2859 N2860 Segment
X2860 N2860 N2861 Segment
X2861 N2861 N2862 Segment
X2862 N2862 N2863 Segment
X2863 N2863 N2864 Segment
X2864 N2864 N2865 Segment
X2865 N2865 N2866 Segment
X2866 N2866 N2867 Segment
X2867 N2867 N2868 Segment
X2868 N2868 N2869 Segment
X2869 N2869 N2870 Segment
X2870 N2870 N2871 Segment
X2871 N2871 N2872 Segment
X2872 N2872 N2873 Segment
X2873 N2873 N2874 Segment
X2874 N2874 N2875 Segment
X2875 N2875 N2876 Segment
X2876 N2876 N2877 Segment
X2877 N2877 N2878 Segment
X2878 N2878 N2879 Segment
X2879 N2879 N2880 Segment
X2880 N2880 N2881 Segment
X2881 N2881 N2882 Segment
X2882 N2882 N2883 Segment
X2883 N2883 N2884 Segment
X2884 N2884 N2885 Segment
X2885 N2885 N2886 Segment
X2886 N2886 N2887 Segment
X2887 N2887 N2888 Segment
X2888 N2888 N2889 Segment
X2889 N2889 N2890 Segment
X2890 N2890 N2891 Segment
X2891 N2891 N2892 Segment
X2892 N2892 N2893 Segment
X2893 N2893 N2894 Segment
X2894 N2894 N2895 Segment
X2895 N2895 N2896 Segment
X2896 N2896 N2897 Segment
X2897 N2897 N2898 Segment
X2898 N2898 N2899 Segment
X2899 N2899 N2900 Segment
X2900 N2900 N2901 Segment
X2901 N2901 N2902 Segment
X2902 N2902 N2903 Segment
X2903 N2903 N2904 Segment
X2904 N2904 N2905 Segment
X2905 N2905 N2906 Segment
X2906 N2906 N2907 Segment
X2907 N2907 N2908 Segment
X2908 N2908 N2909 Segment
X2909 N2909 N2910 Segment
X2910 N2910 N2911 Segment
X2911 N2911 N2912 Segment
X2912 N2912 N2913 Segment
X2913 N2913 N2914 Segment
X2914 N2914 N2915 Segment
X2915 N2915 N2916 Segment
X2916 N2916 N2917 Segment
X2917 N2917 N2918 Segment
X2918 N2918 N2919 Segment
X2919 N2919 N2920 Segment
X2920 N2920 N2921 Segment
X2921 N2921 N2922 Segment
X2922 N2922 N2923 Segment
X2923 N2923 N2924 Segment
X2924 N2924 N2925 Segment
X2925 N2925 N2926 Segment
X2926 N2926 N2927 Segment
X2927 N2927 N2928 Segment
X2928 N2928 N2929 Segment
X2929 N2929 N2930 Segment
X2930 N2930 N2931 Segment
X2931 N2931 N2932 Segment
X2932 N2932 N2933 Segment
X2933 N2933 N2934 Segment
X2934 N2934 N2935 Segment
X2935 N2935 N2936 Segment
X2936 N2936 N2937 Segment
X2937 N2937 N2938 Segment
X2938 N2938 N2939 Segment
X2939 N2939 N2940 Segment
X2940 N2940 N2941 Segment
X2941 N2941 N2942 Segment
X2942 N2942 N2943 Segment
X2943 N2943 N2944 Segment
X2944 N2944 N2945 Segment
X2945 N2945 N2946 Segment
X2946 N2946 N2947 Segment
X2947 N2947 N2948 Segment
X2948 N2948 N2949 Segment
X2949 N2949 N2950 Segment
X2950 N2950 N2951 Segment
X2951 N2951 N2952 Segment
X2952 N2952 N2953 Segment
X2953 N2953 N2954 Segment
X2954 N2954 N2955 Segment
X2955 N2955 N2956 Segment
X2956 N2956 N2957 Segment
X2957 N2957 N2958 Segment
X2958 N2958 N2959 Segment
X2959 N2959 N2960 Segment
X2960 N2960 N2961 Segment
X2961 N2961 N2962 Segment
X2962 N2962 N2963 Segment
X2963 N2963 N2964 Segment
X2964 N2964 N2965 Segment
X2965 N2965 N2966 Segment
X2966 N2966 N2967 Segment
X2967 N2967 N2968 Segment
X2968 N2968 N2969 Segment
X2969 N2969 N2970 Segment
X2970 N2970 N2971 Segment
X2971 N2971 N2972 Segment
X2972 N2972 N2973 Segment
X2973 N2973 N2974 Segment
X2974 N2974 N2975 Segment
X2975 N2975 N2976 Segment
X2976 N2976 N2977 Segment
X2977 N2977 N2978 Segment
X2978 N2978 N2979 Segment
X2979 N2979 N2980 Segment
X2980 N2980 N2981 Segment
X2981 N2981 N2982 Segment
X2982 N2982 N2983 Segment
X2983 N2983 N2984 Segment
X2984 N2984 N2985 Segment
X2985 N2985 N2986 Segment
X2986 N2986 N2987 Segment
X2987 N2987 N2988 Segment
X2988 N2988 N2989 Segment
X2989 N2989 N2990 Segment
X2990 N2990 N2991 Segment
X2991 N2991 N2992 Segment
X2992 N2992 N2993 Segment
X2993 N2993 N2994 Segment
X2994 N2994 N2995 Segment
X2995 N2995 N2996 Segment
X2996 N2996 N2997 Segment
X2997 N2997 N2998 Segment
X2998 N2998 N2999 Segment
X2999 N2999 N3000 Segment
X3000 N3000 N3001 Segment
X3001 N3001 N3002 Segment
X3002 N3002 N3003 Segment
X3003 N3003 N3004 Segment
X3004 N3004 N3005 Segment
X3005 N3005 N3006 Segment
X3006 N3006 N3007 Segment
X3007 N3007 N3008 Segment
X3008 N3008 N3009 Segment
X3009 N3009 N3010 Segment
X3010 N3010 N3011 Segment
X3011 N3011 N3012 Segment
X3012 N3012 N3013 Segment
X3013 N3013 N3014 Segment
X3014 N3014 N3015 Segment
X3015 N3015 N3016 Segment
X3016 N3016 N3017 Segment
X3017 N3017 N3018 Segment
X3018 N3018 N3019 Segment
X3019 N3019 N3020 Segment
X3020 N3020 N3021 Segment
X3021 N3021 N3022 Segment
X3022 N3022 N3023 Segment
X3023 N3023 N3024 Segment
X3024 N3024 N3025 Segment
X3025 N3025 N3026 Segment
X3026 N3026 N3027 Segment
X3027 N3027 N3028 Segment
X3028 N3028 N3029 Segment
X3029 N3029 N3030 Segment
X3030 N3030 N3031 Segment
X3031 N3031 N3032 Segment
X3032 N3032 N3033 Segment
X3033 N3033 N3034 Segment
X3034 N3034 N3035 Segment
X3035 N3035 N3036 Segment
X3036 N3036 N3037 Segment
X3037 N3037 N3038 Segment
X3038 N3038 N3039 Segment
X3039 N3039 N3040 Segment
X3040 N3040 N3041 Segment
X3041 N3041 N3042 Segment
X3042 N3042 N3043 Segment
X3043 N3043 N3044 Segment
X3044 N3044 N3045 Segment
X3045 N3045 N3046 Segment
X3046 N3046 N3047 Segment
X3047 N3047 N3048 Segment
X3048 N3048 N3049 Segment
X3049 N3049 N3050 Segment
X3050 N3050 N3051 Segment
X3051 N3051 N3052 Segment
X3052 N3052 N3053 Segment
X3053 N3053 N3054 Segment
X3054 N3054 N3055 Segment
X3055 N3055 N3056 Segment
X3056 N3056 N3057 Segment
X3057 N3057 N3058 Segment
X3058 N3058 N3059 Segment
X3059 N3059 N3060 Segment
X3060 N3060 N3061 Segment
X3061 N3061 N3062 Segment
X3062 N3062 N3063 Segment
X3063 N3063 N3064 Segment
X3064 N3064 N3065 Segment
X3065 N3065 N3066 Segment
X3066 N3066 N3067 Segment
X3067 N3067 N3068 Segment
X3068 N3068 N3069 Segment
X3069 N3069 N3070 Segment
X3070 N3070 N3071 Segment
X3071 N3071 N3072 Segment
X3072 N3072 N3073 Segment
X3073 N3073 N3074 Segment
X3074 N3074 N3075 Segment
X3075 N3075 N3076 Segment
X3076 N3076 N3077 Segment
X3077 N3077 N3078 Segment
X3078 N3078 N3079 Segment
X3079 N3079 N3080 Segment
X3080 N3080 N3081 Segment
X3081 N3081 N3082 Segment
X3082 N3082 N3083 Segment
X3083 N3083 N3084 Segment
X3084 N3084 N3085 Segment
X3085 N3085 N3086 Segment
X3086 N3086 N3087 Segment
X3087 N3087 N3088 Segment
X3088 N3088 N3089 Segment
X3089 N3089 N3090 Segment
X3090 N3090 N3091 Segment
X3091 N3091 N3092 Segment
X3092 N3092 N3093 Segment
X3093 N3093 N3094 Segment
X3094 N3094 N3095 Segment
X3095 N3095 N3096 Segment
X3096 N3096 N3097 Segment
X3097 N3097 N3098 Segment
X3098 N3098 N3099 Segment
X3099 N3099 N3100 Segment
X3100 N3100 N3101 Segment
X3101 N3101 N3102 Segment
X3102 N3102 N3103 Segment
X3103 N3103 N3104 Segment
X3104 N3104 N3105 Segment
X3105 N3105 N3106 Segment
X3106 N3106 N3107 Segment
X3107 N3107 N3108 Segment
X3108 N3108 N3109 Segment
X3109 N3109 N3110 Segment
X3110 N3110 N3111 Segment
X3111 N3111 N3112 Segment
X3112 N3112 N3113 Segment
X3113 N3113 N3114 Segment
X3114 N3114 N3115 Segment
X3115 N3115 N3116 Segment
X3116 N3116 N3117 Segment
X3117 N3117 N3118 Segment
X3118 N3118 N3119 Segment
X3119 N3119 N3120 Segment
X3120 N3120 N3121 Segment
X3121 N3121 N3122 Segment
X3122 N3122 N3123 Segment
X3123 N3123 N3124 Segment
X3124 N3124 N3125 Segment
X3125 N3125 N3126 Segment
X3126 N3126 N3127 Segment
X3127 N3127 N3128 Segment
X3128 N3128 N3129 Segment
X3129 N3129 N3130 Segment
X3130 N3130 N3131 Segment
X3131 N3131 N3132 Segment
X3132 N3132 N3133 Segment
X3133 N3133 N3134 Segment
X3134 N3134 N3135 Segment
X3135 N3135 N3136 Segment
X3136 N3136 N3137 Segment
X3137 N3137 N3138 Segment
X3138 N3138 N3139 Segment
X3139 N3139 N3140 Segment
X3140 N3140 N3141 Segment
X3141 N3141 N3142 Segment
X3142 N3142 N3143 Segment
X3143 N3143 N3144 Segment
X3144 N3144 N3145 Segment
X3145 N3145 N3146 Segment
X3146 N3146 N3147 Segment
X3147 N3147 N3148 Segment
X3148 N3148 N3149 Segment
X3149 N3149 N3150 Segment
X3150 N3150 N3151 Segment
X3151 N3151 N3152 Segment
X3152 N3152 N3153 Segment
X3153 N3153 N3154 Segment
X3154 N3154 N3155 Segment
X3155 N3155 N3156 Segment
X3156 N3156 N3157 Segment
X3157 N3157 N3158 Segment
X3158 N3158 N3159 Segment
X3159 N3159 N3160 Segment
X3160 N3160 N3161 Segment
X3161 N3161 N3162 Segment
X3162 N3162 N3163 Segment
X3163 N3163 N3164 Segment
X3164 N3164 N3165 Segment
X3165 N3165 N3166 Segment
X3166 N3166 N3167 Segment
X3167 N3167 N3168 Segment
X3168 N3168 N3169 Segment
X3169 N3169 N3170 Segment
X3170 N3170 N3171 Segment
X3171 N3171 N3172 Segment
X3172 N3172 N3173 Segment
X3173 N3173 N3174 Segment
X3174 N3174 N3175 Segment
X3175 N3175 N3176 Segment
X3176 N3176 N3177 Segment
X3177 N3177 N3178 Segment
X3178 N3178 N3179 Segment
X3179 N3179 N3180 Segment
X3180 N3180 N3181 Segment
X3181 N3181 N3182 Segment
X3182 N3182 N3183 Segment
X3183 N3183 N3184 Segment
X3184 N3184 N3185 Segment
X3185 N3185 N3186 Segment
X3186 N3186 N3187 Segment
X3187 N3187 N3188 Segment
X3188 N3188 N3189 Segment
X3189 N3189 N3190 Segment
X3190 N3190 N3191 Segment
X3191 N3191 N3192 Segment
X3192 N3192 N3193 Segment
X3193 N3193 N3194 Segment
X3194 N3194 N3195 Segment
X3195 N3195 N3196 Segment
X3196 N3196 N3197 Segment
X3197 N3197 N3198 Segment
X3198 N3198 N3199 Segment
X3199 N3199 N3200 Segment
X3200 N3200 N3201 Segment
X3201 N3201 N3202 Segment
X3202 N3202 N3203 Segment
X3203 N3203 N3204 Segment
X3204 N3204 N3205 Segment
X3205 N3205 N3206 Segment
X3206 N3206 N3207 Segment
X3207 N3207 N3208 Segment
X3208 N3208 N3209 Segment
X3209 N3209 N3210 Segment
X3210 N3210 N3211 Segment
X3211 N3211 N3212 Segment
X3212 N3212 N3213 Segment
X3213 N3213 N3214 Segment
X3214 N3214 N3215 Segment
X3215 N3215 N3216 Segment
X3216 N3216 N3217 Segment
X3217 N3217 N3218 Segment
X3218 N3218 N3219 Segment
X3219 N3219 N3220 Segment
X3220 N3220 N3221 Segment
X3221 N3221 N3222 Segment
X3222 N3222 N3223 Segment
X3223 N3223 N3224 Segment
X3224 N3224 N3225 Segment
X3225 N3225 N3226 Segment
X3226 N3226 N3227 Segment
X3227 N3227 N3228 Segment
X3228 N3228 N3229 Segment
X3229 N3229 N3230 Segment
X3230 N3230 N3231 Segment
X3231 N3231 N3232 Segment
X3232 N3232 N3233 Segment
X3233 N3233 N3234 Segment
X3234 N3234 N3235 Segment
X3235 N3235 N3236 Segment
X3236 N3236 N3237 Segment
X3237 N3237 N3238 Segment
X3238 N3238 N3239 Segment
X3239 N3239 N3240 Segment
X3240 N3240 N3241 Segment
X3241 N3241 N3242 Segment
X3242 N3242 N3243 Segment
X3243 N3243 N3244 Segment
X3244 N3244 N3245 Segment
X3245 N3245 N3246 Segment
X3246 N3246 N3247 Segment
X3247 N3247 N3248 Segment
X3248 N3248 N3249 Segment
X3249 N3249 N3250 Segment
X3250 N3250 N3251 Segment
X3251 N3251 N3252 Segment
X3252 N3252 N3253 Segment
X3253 N3253 N3254 Segment
X3254 N3254 N3255 Segment
X3255 N3255 N3256 Segment
X3256 N3256 N3257 Segment
X3257 N3257 N3258 Segment
X3258 N3258 N3259 Segment
X3259 N3259 N3260 Segment
X3260 N3260 N3261 Segment
X3261 N3261 N3262 Segment
X3262 N3262 N3263 Segment
X3263 N3263 N3264 Segment
X3264 N3264 N3265 Segment
X3265 N3265 N3266 Segment
X3266 N3266 N3267 Segment
X3267 N3267 N3268 Segment
X3268 N3268 N3269 Segment
X3269 N3269 N3270 Segment
X3270 N3270 N3271 Segment
X3271 N3271 N3272 Segment
X3272 N3272 N3273 Segment
X3273 N3273 N3274 Segment
X3274 N3274 N3275 Segment
X3275 N3275 N3276 Segment
X3276 N3276 N3277 Segment
X3277 N3277 N3278 Segment
X3278 N3278 N3279 Segment
X3279 N3279 N3280 Segment
X3280 N3280 N3281 Segment
X3281 N3281 N3282 Segment
X3282 N3282 N3283 Segment
X3283 N3283 N3284 Segment
X3284 N3284 N3285 Segment
X3285 N3285 N3286 Segment
X3286 N3286 N3287 Segment
X3287 N3287 N3288 Segment
X3288 N3288 N3289 Segment
X3289 N3289 N3290 Segment
X3290 N3290 N3291 Segment
X3291 N3291 N3292 Segment
X3292 N3292 N3293 Segment
X3293 N3293 N3294 Segment
X3294 N3294 N3295 Segment
X3295 N3295 N3296 Segment
X3296 N3296 N3297 Segment
X3297 N3297 N3298 Segment
X3298 N3298 N3299 Segment
X3299 N3299 N3300 Segment
X3300 N3300 N3301 Segment
X3301 N3301 N3302 Segment
X3302 N3302 N3303 Segment
X3303 N3303 N3304 Segment
X3304 N3304 N3305 Segment
X3305 N3305 N3306 Segment
X3306 N3306 N3307 Segment
X3307 N3307 N3308 Segment
X3308 N3308 N3309 Segment
X3309 N3309 N3310 Segment
X3310 N3310 N3311 Segment
X3311 N3311 N3312 Segment
X3312 N3312 N3313 Segment
X3313 N3313 N3314 Segment
X3314 N3314 N3315 Segment
X3315 N3315 N3316 Segment
X3316 N3316 N3317 Segment
X3317 N3317 N3318 Segment
X3318 N3318 N3319 Segment
X3319 N3319 N3320 Segment
X3320 N3320 N3321 Segment
X3321 N3321 N3322 Segment
X3322 N3322 N3323 Segment
X3323 N3323 N3324 Segment
X3324 N3324 N3325 Segment
X3325 N3325 N3326 Segment
X3326 N3326 N3327 Segment
X3327 N3327 N3328 Segment
X3328 N3328 N3329 Segment
X3329 N3329 N3330 Segment
X3330 N3330 N3331 Segment
X3331 N3331 N3332 Segment
X3332 N3332 N3333 Segment
X3333 N3333 N3334 Segment
X3334 N3334 N3335 Segment
X3335 N3335 N3336 Segment
X3336 N3336 N3337 Segment
X3337 N3337 N3338 Segment
X3338 N3338 N3339 Segment
X3339 N3339 N3340 Segment
X3340 N3340 N3341 Segment
X3341 N3341 N3342 Segment
X3342 N3342 N3343 Segment
X3343 N3343 N3344 Segment
X3344 N3344 N3345 Segment
X3345 N3345 N3346 Segment
X3346 N3346 N3347 Segment
X3347 N3347 N3348 Segment
X3348 N3348 N3349 Segment
X3349 N3349 N3350 Segment
X3350 N3350 N3351 Segment
X3351 N3351 N3352 Segment
X3352 N3352 N3353 Segment
X3353 N3353 N3354 Segment
X3354 N3354 N3355 Segment
X3355 N3355 N3356 Segment
X3356 N3356 N3357 Segment
X3357 N3357 N3358 Segment
X3358 N3358 N3359 Segment
X3359 N3359 N3360 Segment
X3360 N3360 N3361 Segment
X3361 N3361 N3362 Segment
X3362 N3362 N3363 Segment
X3363 N3363 N3364 Segment
X3364 N3364 N3365 Segment
X3365 N3365 N3366 Segment
X3366 N3366 N3367 Segment
X3367 N3367 N3368 Segment
X3368 N3368 N3369 Segment
X3369 N3369 N3370 Segment
X3370 N3370 N3371 Segment
X3371 N3371 N3372 Segment
X3372 N3372 N3373 Segment
X3373 N3373 N3374 Segment
X3374 N3374 N3375 Segment
X3375 N3375 N3376 Segment
X3376 N3376 N3377 Segment
X3377 N3377 N3378 Segment
X3378 N3378 N3379 Segment
X3379 N3379 N3380 Segment
X3380 N3380 N3381 Segment
X3381 N3381 N3382 Segment
X3382 N3382 N3383 Segment
X3383 N3383 N3384 Segment
X3384 N3384 N3385 Segment
X3385 N3385 N3386 Segment
X3386 N3386 N3387 Segment
X3387 N3387 N3388 Segment
X3388 N3388 N3389 Segment
X3389 N3389 N3390 Segment
X3390 N3390 N3391 Segment
X3391 N3391 N3392 Segment
X3392 N3392 N3393 Segment
X3393 N3393 N3394 Segment
X3394 N3394 N3395 Segment
X3395 N3395 N3396 Segment
X3396 N3396 N3397 Segment
X3397 N3397 N3398 Segment
X3398 N3398 N3399 Segment
X3399 N3399 N3400 Segment
X3400 N3400 N3401 Segment
X3401 N3401 N3402 Segment
X3402 N3402 N3403 Segment
X3403 N3403 N3404 Segment
X3404 N3404 N3405 Segment
X3405 N3405 N3406 Segment
X3406 N3406 N3407 Segment
X3407 N3407 N3408 Segment
X3408 N3408 N3409 Segment
X3409 N3409 N3410 Segment
X3410 N3410 N3411 Segment
X3411 N3411 N3412 Segment
X3412 N3412 N3413 Segment
X3413 N3413 N3414 Segment
X3414 N3414 N3415 Segment
X3415 N3415 N3416 Segment
X3416 N3416 N3417 Segment
X3417 N3417 N3418 Segment
X3418 N3418 N3419 Segment
X3419 N3419 N3420 Segment
X3420 N3420 N3421 Segment
X3421 N3421 N3422 Segment
X3422 N3422 N3423 Segment
X3423 N3423 N3424 Segment
X3424 N3424 N3425 Segment
X3425 N3425 N3426 Segment
X3426 N3426 N3427 Segment
X3427 N3427 N3428 Segment
X3428 N3428 N3429 Segment
X3429 N3429 N3430 Segment
X3430 N3430 N3431 Segment
X3431 N3431 N3432 Segment
X3432 N3432 N3433 Segment
X3433 N3433 N3434 Segment
X3434 N3434 N3435 Segment
X3435 N3435 N3436 Segment
X3436 N3436 N3437 Segment
X3437 N3437 N3438 Segment
X3438 N3438 N3439 Segment
X3439 N3439 N3440 Segment
X3440 N3440 N3441 Segment
X3441 N3441 N3442 Segment
X3442 N3442 N3443 Segment
X3443 N3443 N3444 Segment
X3444 N3444 N3445 Segment
X3445 N3445 N3446 Segment
X3446 N3446 N3447 Segment
X3447 N3447 N3448 Segment
X3448 N3448 N3449 Segment
X3449 N3449 N3450 Segment
X3450 N3450 N3451 Segment
X3451 N3451 N3452 Segment
X3452 N3452 N3453 Segment
X3453 N3453 N3454 Segment
X3454 N3454 N3455 Segment
X3455 N3455 N3456 Segment
X3456 N3456 N3457 Segment
X3457 N3457 N3458 Segment
X3458 N3458 N3459 Segment
X3459 N3459 N3460 Segment
X3460 N3460 N3461 Segment
X3461 N3461 N3462 Segment
X3462 N3462 N3463 Segment
X3463 N3463 N3464 Segment
X3464 N3464 N3465 Segment
X3465 N3465 N3466 Segment
X3466 N3466 N3467 Segment
X3467 N3467 N3468 Segment
X3468 N3468 N3469 Segment
X3469 N3469 N3470 Segment
X3470 N3470 N3471 Segment
X3471 N3471 N3472 Segment
X3472 N3472 N3473 Segment
X3473 N3473 N3474 Segment
X3474 N3474 N3475 Segment
X3475 N3475 N3476 Segment
X3476 N3476 N3477 Segment
X3477 N3477 N3478 Segment
X3478 N3478 N3479 Segment
X3479 N3479 N3480 Segment
X3480 N3480 N3481 Segment
X3481 N3481 N3482 Segment
X3482 N3482 N3483 Segment
X3483 N3483 N3484 Segment
X3484 N3484 N3485 Segment
X3485 N3485 N3486 Segment
X3486 N3486 N3487 Segment
X3487 N3487 N3488 Segment
X3488 N3488 N3489 Segment
X3489 N3489 N3490 Segment
X3490 N3490 N3491 Segment
X3491 N3491 N3492 Segment
X3492 N3492 N3493 Segment
X3493 N3493 N3494 Segment
X3494 N3494 N3495 Segment
X3495 N3495 N3496 Segment
X3496 N3496 N3497 Segment
X3497 N3497 N3498 Segment
X3498 N3498 N3499 Segment
X3499 N3499 N3500 Segment
X3500 N3500 N3501 Segment
X3501 N3501 N3502 Segment
X3502 N3502 N3503 Segment
X3503 N3503 N3504 Segment
X3504 N3504 N3505 Segment
X3505 N3505 N3506 Segment
X3506 N3506 N3507 Segment
X3507 N3507 N3508 Segment
X3508 N3508 N3509 Segment
X3509 N3509 N3510 Segment
X3510 N3510 N3511 Segment
X3511 N3511 N3512 Segment
X3512 N3512 N3513 Segment
X3513 N3513 N3514 Segment
X3514 N3514 N3515 Segment
X3515 N3515 N3516 Segment
X3516 N3516 N3517 Segment
X3517 N3517 N3518 Segment
X3518 N3518 N3519 Segment
X3519 N3519 N3520 Segment
X3520 N3520 N3521 Segment
X3521 N3521 N3522 Segment
X3522 N3522 N3523 Segment
X3523 N3523 N3524 Segment
X3524 N3524 N3525 Segment
X3525 N3525 N3526 Segment
X3526 N3526 N3527 Segment
X3527 N3527 N3528 Segment
X3528 N3528 N3529 Segment
X3529 N3529 N3530 Segment
X3530 N3530 N3531 Segment
X3531 N3531 N3532 Segment
X3532 N3532 N3533 Segment
X3533 N3533 N3534 Segment
X3534 N3534 N3535 Segment
X3535 N3535 N3536 Segment
X3536 N3536 N3537 Segment
X3537 N3537 N3538 Segment
X3538 N3538 N3539 Segment
X3539 N3539 N3540 Segment
X3540 N3540 N3541 Segment
X3541 N3541 N3542 Segment
X3542 N3542 N3543 Segment
X3543 N3543 N3544 Segment
X3544 N3544 N3545 Segment
X3545 N3545 N3546 Segment
X3546 N3546 N3547 Segment
X3547 N3547 N3548 Segment
X3548 N3548 N3549 Segment
X3549 N3549 N3550 Segment
X3550 N3550 N3551 Segment
X3551 N3551 N3552 Segment
X3552 N3552 N3553 Segment
X3553 N3553 N3554 Segment
X3554 N3554 N3555 Segment
X3555 N3555 N3556 Segment
X3556 N3556 N3557 Segment
X3557 N3557 N3558 Segment
X3558 N3558 N3559 Segment
X3559 N3559 N3560 Segment
X3560 N3560 N3561 Segment
X3561 N3561 N3562 Segment
X3562 N3562 N3563 Segment
X3563 N3563 N3564 Segment
X3564 N3564 N3565 Segment
X3565 N3565 N3566 Segment
X3566 N3566 N3567 Segment
X3567 N3567 N3568 Segment
X3568 N3568 N3569 Segment
X3569 N3569 N3570 Segment
X3570 N3570 N3571 Segment
X3571 N3571 N3572 Segment
X3572 N3572 N3573 Segment
X3573 N3573 N3574 Segment
X3574 N3574 N3575 Segment
X3575 N3575 N3576 Segment
X3576 N3576 N3577 Segment
X3577 N3577 N3578 Segment
X3578 N3578 N3579 Segment
X3579 N3579 N3580 Segment
X3580 N3580 N3581 Segment
X3581 N3581 N3582 Segment
X3582 N3582 N3583 Segment
X3583 N3583 N3584 Segment
X3584 N3584 N3585 Segment
X3585 N3585 N3586 Segment
X3586 N3586 N3587 Segment
X3587 N3587 N3588 Segment
X3588 N3588 N3589 Segment
X3589 N3589 N3590 Segment
X3590 N3590 N3591 Segment
X3591 N3591 N3592 Segment
X3592 N3592 N3593 Segment
X3593 N3593 N3594 Segment
X3594 N3594 N3595 Segment
X3595 N3595 N3596 Segment
X3596 N3596 N3597 Segment
X3597 N3597 N3598 Segment
X3598 N3598 N3599 Segment
X3599 N3599 N3600 Segment
X3600 N3600 N3601 Segment
X3601 N3601 N3602 Segment
X3602 N3602 N3603 Segment
X3603 N3603 N3604 Segment
X3604 N3604 N3605 Segment
X3605 N3605 N3606 Segment
X3606 N3606 N3607 Segment
X3607 N3607 N3608 Segment
X3608 N3608 N3609 Segment
X3609 N3609 N3610 Segment
X3610 N3610 N3611 Segment
X3611 N3611 N3612 Segment
X3612 N3612 N3613 Segment
X3613 N3613 N3614 Segment
X3614 N3614 N3615 Segment
X3615 N3615 N3616 Segment
X3616 N3616 N3617 Segment
X3617 N3617 N3618 Segment
X3618 N3618 N3619 Segment
X3619 N3619 N3620 Segment
X3620 N3620 N3621 Segment
X3621 N3621 N3622 Segment
X3622 N3622 N3623 Segment
X3623 N3623 N3624 Segment
X3624 N3624 N3625 Segment
X3625 N3625 N3626 Segment
X3626 N3626 N3627 Segment
X3627 N3627 N3628 Segment
X3628 N3628 N3629 Segment
X3629 N3629 N3630 Segment
X3630 N3630 N3631 Segment
X3631 N3631 N3632 Segment
X3632 N3632 N3633 Segment
X3633 N3633 N3634 Segment
X3634 N3634 N3635 Segment
X3635 N3635 N3636 Segment
X3636 N3636 N3637 Segment
X3637 N3637 N3638 Segment
X3638 N3638 N3639 Segment
X3639 N3639 N3640 Segment
X3640 N3640 N3641 Segment
X3641 N3641 N3642 Segment
X3642 N3642 N3643 Segment
X3643 N3643 N3644 Segment
X3644 N3644 N3645 Segment
X3645 N3645 N3646 Segment
X3646 N3646 N3647 Segment
X3647 N3647 N3648 Segment
X3648 N3648 N3649 Segment
X3649 N3649 N3650 Segment
X3650 N3650 N3651 Segment
X3651 N3651 N3652 Segment
X3652 N3652 N3653 Segment
X3653 N3653 N3654 Segment
X3654 N3654 N3655 Segment
X3655 N3655 N3656 Segment
X3656 N3656 N3657 Segment
X3657 N3657 N3658 Segment
X3658 N3658 N3659 Segment
X3659 N3659 N3660 Segment
X3660 N3660 N3661 Segment
X3661 N3661 N3662 Segment
X3662 N3662 N3663 Segment
X3663 N3663 N3664 Segment
X3664 N3664 N3665 Segment
X3665 N3665 N3666 Segment
X3666 N3666 N3667 Segment
X3667 N3667 N3668 Segment
X3668 N3668 N3669 Segment
X3669 N3669 N3670 Segment
X3670 N3670 N3671 Segment
X3671 N3671 N3672 Segment
X3672 N3672 N3673 Segment
X3673 N3673 N3674 Segment
X3674 N3674 N3675 Segment
X3675 N3675 N3676 Segment
X3676 N3676 N3677 Segment
X3677 N3677 N3678 Segment
X3678 N3678 N3679 Segment
X3679 N3679 N3680 Segment
X3680 N3680 N3681 Segment
X3681 N3681 N3682 Segment
X3682 N3682 N3683 Segment
X3683 N3683 N3684 Segment
X3684 N3684 N3685 Segment
X3685 N3685 N3686 Segment
X3686 N3686 N3687 Segment
X3687 N3687 N3688 Segment
X3688 N3688 N3689 Segment
X3689 N3689 N3690 Segment
X3690 N3690 N3691 Segment
X3691 N3691 N3692 Segment
X3692 N3692 N3693 Segment
X3693 N3693 N3694 Segment
X3694 N3694 N3695 Segment
X3695 N3695 N3696 Segment
X3696 N3696 N3697 Segment
X3697 N3697 N3698 Segment
X3698 N3698 N3699 Segment
X3699 N3699 N3700 Segment
X3700 N3700 N3701 Segment
X3701 N3701 N3702 Segment
X3702 N3702 N3703 Segment
X3703 N3703 N3704 Segment
X3704 N3704 N3705 Segment
X3705 N3705 N3706 Segment
X3706 N3706 N3707 Segment
X3707 N3707 N3708 Segment
X3708 N3708 N3709 Segment
X3709 N3709 N3710 Segment
X3710 N3710 N3711 Segment
X3711 N3711 N3712 Segment
X3712 N3712 N3713 Segment
X3713 N3713 N3714 Segment
X3714 N3714 N3715 Segment
X3715 N3715 N3716 Segment
X3716 N3716 N3717 Segment
X3717 N3717 N3718 Segment
X3718 N3718 N3719 Segment
X3719 N3719 N3720 Segment
X3720 N3720 N3721 Segment
X3721 N3721 N3722 Segment
X3722 N3722 N3723 Segment
X3723 N3723 N3724 Segment
X3724 N3724 N3725 Segment
X3725 N3725 N3726 Segment
X3726 N3726 N3727 Segment
X3727 N3727 N3728 Segment
X3728 N3728 N3729 Segment
X3729 N3729 N3730 Segment
X3730 N3730 N3731 Segment
X3731 N3731 N3732 Segment
X3732 N3732 N3733 Segment
X3733 N3733 N3734 Segment
X3734 N3734 N3735 Segment
X3735 N3735 N3736 Segment
X3736 N3736 N3737 Segment
X3737 N3737 N3738 Segment
X3738 N3738 N3739 Segment
X3739 N3739 N3740 Segment
X3740 N3740 N3741 Segment
X3741 N3741 N3742 Segment
X3742 N3742 N3743 Segment
X3743 N3743 N3744 Segment
X3744 N3744 N3745 Segment
X3745 N3745 N3746 Segment
X3746 N3746 N3747 Segment
X3747 N3747 N3748 Segment
X3748 N3748 N3749 Segment
X3749 N3749 N3750 Segment
X3750 N3750 N3751 Segment
X3751 N3751 N3752 Segment
X3752 N3752 N3753 Segment
X3753 N3753 N3754 Segment
X3754 N3754 N3755 Segment
X3755 N3755 N3756 Segment
X3756 N3756 N3757 Segment
X3757 N3757 N3758 Segment
X3758 N3758 N3759 Segment
X3759 N3759 N3760 Segment
X3760 N3760 N3761 Segment
X3761 N3761 N3762 Segment
X3762 N3762 N3763 Segment
X3763 N3763 N3764 Segment
X3764 N3764 N3765 Segment
X3765 N3765 N3766 Segment
X3766 N3766 N3767 Segment
X3767 N3767 N3768 Segment
X3768 N3768 N3769 Segment
X3769 N3769 N3770 Segment
X3770 N3770 N3771 Segment
X3771 N3771 N3772 Segment
X3772 N3772 N3773 Segment
X3773 N3773 N3774 Segment
X3774 N3774 N3775 Segment
X3775 N3775 N3776 Segment
X3776 N3776 N3777 Segment
X3777 N3777 N3778 Segment
X3778 N3778 N3779 Segment
X3779 N3779 N3780 Segment
X3780 N3780 N3781 Segment
X3781 N3781 N3782 Segment
X3782 N3782 N3783 Segment
X3783 N3783 N3784 Segment
X3784 N3784 N3785 Segment
X3785 N3785 N3786 Segment
X3786 N3786 N3787 Segment
X3787 N3787 N3788 Segment
X3788 N3788 N3789 Segment
X3789 N3789 N3790 Segment
X3790 N3790 N3791 Segment
X3791 N3791 N3792 Segment
X3792 N3792 N3793 Segment
X3793 N3793 N3794 Segment
X3794 N3794 N3795 Segment
X3795 N3795 N3796 Segment
X3796 N3796 N3797 Segment
X3797 N3797 N3798 Segment
X3798 N3798 N3799 Segment
X3799 N3799 N3800 Segment
X3800 N3800 N3801 Segment
X3801 N3801 N3802 Segment
X3802 N3802 N3803 Segment
X3803 N3803 N3804 Segment
X3804 N3804 N3805 Segment
X3805 N3805 N3806 Segment
X3806 N3806 N3807 Segment
X3807 N3807 N3808 Segment
X3808 N3808 N3809 Segment
X3809 N3809 N3810 Segment
X3810 N3810 N3811 Segment
X3811 N3811 N3812 Segment
X3812 N3812 N3813 Segment
X3813 N3813 N3814 Segment
X3814 N3814 N3815 Segment
X3815 N3815 N3816 Segment
X3816 N3816 N3817 Segment
X3817 N3817 N3818 Segment
X3818 N3818 N3819 Segment
X3819 N3819 N3820 Segment
X3820 N3820 N3821 Segment
X3821 N3821 N3822 Segment
X3822 N3822 N3823 Segment
X3823 N3823 N3824 Segment
X3824 N3824 N3825 Segment
X3825 N3825 N3826 Segment
X3826 N3826 N3827 Segment
X3827 N3827 N3828 Segment
X3828 N3828 N3829 Segment
X3829 N3829 N3830 Segment
X3830 N3830 N3831 Segment
X3831 N3831 N3832 Segment
X3832 N3832 N3833 Segment
X3833 N3833 N3834 Segment
X3834 N3834 N3835 Segment
X3835 N3835 N3836 Segment
X3836 N3836 N3837 Segment
X3837 N3837 N3838 Segment
X3838 N3838 N3839 Segment
X3839 N3839 N3840 Segment
X3840 N3840 N3841 Segment
X3841 N3841 N3842 Segment
X3842 N3842 N3843 Segment
X3843 N3843 N3844 Segment
X3844 N3844 N3845 Segment
X3845 N3845 N3846 Segment
X3846 N3846 N3847 Segment
X3847 N3847 N3848 Segment
X3848 N3848 N3849 Segment
X3849 N3849 N3850 Segment
X3850 N3850 N3851 Segment
X3851 N3851 N3852 Segment
X3852 N3852 N3853 Segment
X3853 N3853 N3854 Segment
X3854 N3854 N3855 Segment
X3855 N3855 N3856 Segment
X3856 N3856 N3857 Segment
X3857 N3857 N3858 Segment
X3858 N3858 N3859 Segment
X3859 N3859 N3860 Segment
X3860 N3860 N3861 Segment
X3861 N3861 N3862 Segment
X3862 N3862 N3863 Segment
X3863 N3863 N3864 Segment
X3864 N3864 N3865 Segment
X3865 N3865 N3866 Segment
X3866 N3866 N3867 Segment
X3867 N3867 N3868 Segment
X3868 N3868 N3869 Segment
X3869 N3869 N3870 Segment
X3870 N3870 N3871 Segment
X3871 N3871 N3872 Segment
X3872 N3872 N3873 Segment
X3873 N3873 N3874 Segment
X3874 N3874 N3875 Segment
X3875 N3875 N3876 Segment
X3876 N3876 N3877 Segment
X3877 N3877 N3878 Segment
X3878 N3878 N3879 Segment
X3879 N3879 N3880 Segment
X3880 N3880 N3881 Segment
X3881 N3881 N3882 Segment
X3882 N3882 N3883 Segment
X3883 N3883 N3884 Segment
X3884 N3884 N3885 Segment
X3885 N3885 N3886 Segment
X3886 N3886 N3887 Segment
X3887 N3887 N3888 Segment
X3888 N3888 N3889 Segment
X3889 N3889 N3890 Segment
X3890 N3890 N3891 Segment
X3891 N3891 N3892 Segment
X3892 N3892 N3893 Segment
X3893 N3893 N3894 Segment
X3894 N3894 N3895 Segment
X3895 N3895 N3896 Segment
X3896 N3896 N3897 Segment
X3897 N3897 N3898 Segment
X3898 N3898 N3899 Segment
X3899 N3899 N3900 Segment
X3900 N3900 N3901 Segment
X3901 N3901 N3902 Segment
X3902 N3902 N3903 Segment
X3903 N3903 N3904 Segment
X3904 N3904 N3905 Segment
X3905 N3905 N3906 Segment
X3906 N3906 N3907 Segment
X3907 N3907 N3908 Segment
X3908 N3908 N3909 Segment
X3909 N3909 N3910 Segment
X3910 N3910 N3911 Segment
X3911 N3911 N3912 Segment
X3912 N3912 N3913 Segment
X3913 N3913 N3914 Segment
X3914 N3914 N3915 Segment
X3915 N3915 N3916 Segment
X3916 N3916 N3917 Segment
X3917 N3917 N3918 Segment
X3918 N3918 N3919 Segment
X3919 N3919 N3920 Segment
X3920 N3920 N3921 Segment
X3921 N3921 N3922 Segment
X3922 N3922 N3923 Segment
X3923 N3923 N3924 Segment
X3924 N3924 N3925 Segment
X3925 N3925 N3926 Segment
X3926 N3926 N3927 Segment
X3927 N3927 N3928 Segment
X3928 N3928 N3929 Segment
X3929 N3929 N3930 Segment
X3930 N3930 N3931 Segment
X3931 N3931 N3932 Segment
X3932 N3932 N3933 Segment
X3933 N3933 N3934 Segment
X3934 N3934 N3935 Segment
X3935 N3935 N3936 Segment
X3936 N3936 N3937 Segment
X3937 N3937 N3938 Segment
X3938 N3938 N3939 Segment
X3939 N3939 N3940 Segment
X3940 N3940 N3941 Segment
X3941 N3941 N3942 Segment
X3942 N3942 N3943 Segment
X3943 N3943 N3944 Segment
X3944 N3944 N3945 Segment
X3945 N3945 N3946 Segment
X3946 N3946 N3947 Segment
X3947 N3947 N3948 Segment
X3948 N3948 N3949 Segment
X3949 N3949 N3950 Segment
X3950 N3950 N3951 Segment
X3951 N3951 N3952 Segment
X3952 N3952 N3953 Segment
X3953 N3953 N3954 Segment
X3954 N3954 N3955 Segment
X3955 N3955 N3956 Segment
X3956 N3956 N3957 Segment
X3957 N3957 N3958 Segment
X3958 N3958 N3959 Segment
X3959 N3959 N3960 Segment
X3960 N3960 N3961 Segment
X3961 N3961 N3962 Segment
X3962 N3962 N3963 Segment
X3963 N3963 N3964 Segment
X3964 N3964 N3965 Segment
X3965 N3965 N3966 Segment
X3966 N3966 N3967 Segment
X3967 N3967 N3968 Segment
X3968 N3968 N3969 Segment
X3969 N3969 N3970 Segment
X3970 N3970 N3971 Segment
X3971 N3971 N3972 Segment
X3972 N3972 N3973 Segment
X3973 N3973 N3974 Segment
X3974 N3974 N3975 Segment
X3975 N3975 N3976 Segment
X3976 N3976 N3977 Segment
X3977 N3977 N3978 Segment
X3978 N3978 N3979 Segment
X3979 N3979 N3980 Segment
X3980 N3980 N3981 Segment
X3981 N3981 N3982 Segment
X3982 N3982 N3983 Segment
X3983 N3983 N3984 Segment
X3984 N3984 N3985 Segment
X3985 N3985 N3986 Segment
X3986 N3986 N3987 Segment
X3987 N3987 N3988 Segment
X3988 N3988 N3989 Segment
X3989 N3989 N3990 Segment
X3990 N3990 N3991 Segment
X3991 N3991 N3992 Segment
X3992 N3992 N3993 Segment
X3993 N3993 N3994 Segment
X3994 N3994 N3995 Segment
X3995 N3995 N3996 Segment
X3996 N3996 N3997 Segment
X3997 N3997 N3998 Segment
X3998 N3998 N3999 Segment
X3999 N3999 N4000 Segment
X4000 N4000 N4001 Segment
X4001 N4001 N4002 Segment
X4002 N4002 N4003 Segment
X4003 N4003 N4004 Segment
X4004 N4004 N4005 Segment
X4005 N4005 N4006 Segment
X4006 N4006 N4007 Segment
X4007 N4007 N4008 Segment
X4008 N4008 N4009 Segment
X4009 N4009 N4010 Segment
X4010 N4010 N4011 Segment
X4011 N4011 N4012 Segment
X4012 N4012 N4013 Segment
X4013 N4013 N4014 Segment
X4014 N4014 N4015 Segment
X4015 N4015 N4016 Segment
X4016 N4016 N4017 Segment
X4017 N4017 N4018 Segment
X4018 N4018 N4019 Segment
X4019 N4019 N4020 Segment
X4020 N4020 N4021 Segment
X4021 N4021 N4022 Segment
X4022 N4022 N4023 Segment
X4023 N4023 N4024 Segment
X4024 N4024 N4025 Segment
X4025 N4025 N4026 Segment
X4026 N4026 N4027 Segment
X4027 N4027 N4028 Segment
X4028 N4028 N4029 Segment
X4029 N4029 N4030 Segment
X4030 N4030 N4031 Segment
X4031 N4031 N4032 Segment
X4032 N4032 N4033 Segment
X4033 N4033 N4034 Segment
X4034 N4034 N4035 Segment
X4035 N4035 N4036 Segment
X4036 N4036 N4037 Segment
X4037 N4037 N4038 Segment
X4038 N4038 N4039 Segment
X4039 N4039 N4040 Segment
X4040 N4040 N4041 Segment
X4041 N4041 N4042 Segment
X4042 N4042 N4043 Segment
X4043 N4043 N4044 Segment
X4044 N4044 N4045 Segment
X4045 N4045 N4046 Segment
X4046 N4046 N4047 Segment
X4047 N4047 N4048 Segment
X4048 N4048 N4049 Segment
X4049 N4049 N4050 Segment
X4050 N4050 N4051 Segment
X4051 N4051 N4052 Segment
X4052 N4052 N4053 Segment
X4053 N4053 N4054 Segment
X4054 N4054 N4055 Segment
X4055 N4055 N4056 Segment
X4056 N4056 N4057 Segment
X4057 N4057 N4058 Segment
X4058 N4058 N4059 Segment
X4059 N4059 N4060 Segment
X4060 N4060 N4061 Segment
X4061 N4061 N4062 Segment
X4062 N4062 N4063 Segment
X4063 N4063 N4064 Segment
X4064 N4064 N4065 Segment
X4065 N4065 N4066 Segment
X4066 N4066 N4067 Segment
X4067 N4067 N4068 Segment
X4068 N4068 N4069 Segment
X4069 N4069 N4070 Segment
X4070 N4070 N4071 Segment
X4071 N4071 N4072 Segment
X4072 N4072 N4073 Segment
X4073 N4073 N4074 Segment
X4074 N4074 N4075 Segment
X4075 N4075 N4076 Segment
X4076 N4076 N4077 Segment
X4077 N4077 N4078 Segment
X4078 N4078 N4079 Segment
X4079 N4079 N4080 Segment
X4080 N4080 N4081 Segment
X4081 N4081 N4082 Segment
X4082 N4082 N4083 Segment
X4083 N4083 N4084 Segment
X4084 N4084 N4085 Segment
X4085 N4085 N4086 Segment
X4086 N4086 N4087 Segment
X4087 N4087 N4088 Segment
X4088 N4088 N4089 Segment
X4089 N4089 N4090 Segment
X4090 N4090 N4091 Segment
X4091 N4091 N4092 Segment
X4092 N4092 N4093 Segment
X4093 N4093 N4094 Segment
X4094 N4094 N4095 Segment
X4095 N4095 N4096 Segment
X4096 N4096 N4097 Segment
X4097 N4097 N4098 Segment
X4098 N4098 N4099 Segment
X4099 N4099 N4100 Segment
X4100 N4100 N4101 Segment
X4101 N4101 N4102 Segment
X4102 N4102 N4103 Segment
X4103 N4103 N4104 Segment
X4104 N4104 N4105 Segment
X4105 N4105 N4106 Segment
X4106 N4106 N4107 Segment
X4107 N4107 N4108 Segment
X4108 N4108 N4109 Segment
X4109 N4109 N4110 Segment
X4110 N4110 N4111 Segment
X4111 N4111 N4112 Segment
X4112 N4112 N4113 Segment
X4113 N4113 N4114 Segment
X4114 N4114 N4115 Segment
X4115 N4115 N4116 Segment
X4116 N4116 N4117 Segment
X4117 N4117 N4118 Segment
X4118 N4118 N4119 Segment
X4119 N4119 N4120 Segment
X4120 N4120 N4121 Segment
X4121 N4121 N4122 Segment
X4122 N4122 N4123 Segment
X4123 N4123 N4124 Segment
X4124 N4124 N4125 Segment
X4125 N4125 N4126 Segment
X4126 N4126 N4127 Segment
X4127 N4127 N4128 Segment
X4128 N4128 N4129 Segment
X4129 N4129 N4130 Segment
X4130 N4130 N4131 Segment
X4131 N4131 N4132 Segment
X4132 N4132 N4133 Segment
X4133 N4133 N4134 Segment
X4134 N4134 N4135 Segment
X4135 N4135 N4136 Segment
X4136 N4136 N4137 Segment
X4137 N4137 N4138 Segment
X4138 N4138 N4139 Segment
X4139 N4139 N4140 Segment
X4140 N4140 N4141 Segment
X4141 N4141 N4142 Segment
X4142 N4142 N4143 Segment
X4143 N4143 N4144 Segment
X4144 N4144 N4145 Segment
X4145 N4145 N4146 Segment
X4146 N4146 N4147 Segment
X4147 N4147 N4148 Segment
X4148 N4148 N4149 Segment
X4149 N4149 N4150 Segment
X4150 N4150 N4151 Segment
X4151 N4151 N4152 Segment
X4152 N4152 N4153 Segment
X4153 N4153 N4154 Segment
X4154 N4154 N4155 Segment
X4155 N4155 N4156 Segment
X4156 N4156 N4157 Segment
X4157 N4157 N4158 Segment
X4158 N4158 N4159 Segment
X4159 N4159 N4160 Segment
X4160 N4160 N4161 Segment
X4161 N4161 N4162 Segment
X4162 N4162 N4163 Segment
X4163 N4163 N4164 Segment
X4164 N4164 N4165 Segment
X4165 N4165 N4166 Segment
X4166 N4166 N4167 Segment
X4167 N4167 N4168 Segment
X4168 N4168 N4169 Segment
X4169 N4169 N4170 Segment
X4170 N4170 N4171 Segment
X4171 N4171 N4172 Segment
X4172 N4172 N4173 Segment
X4173 N4173 N4174 Segment
X4174 N4174 N4175 Segment
X4175 N4175 N4176 Segment
X4176 N4176 N4177 Segment
X4177 N4177 N4178 Segment
X4178 N4178 N4179 Segment
X4179 N4179 N4180 Segment
X4180 N4180 N4181 Segment
X4181 N4181 N4182 Segment
X4182 N4182 N4183 Segment
X4183 N4183 N4184 Segment
X4184 N4184 N4185 Segment
X4185 N4185 N4186 Segment
X4186 N4186 N4187 Segment
X4187 N4187 N4188 Segment
X4188 N4188 N4189 Segment
X4189 N4189 N4190 Segment
X4190 N4190 N4191 Segment
X4191 N4191 N4192 Segment
X4192 N4192 N4193 Segment
X4193 N4193 N4194 Segment
X4194 N4194 N4195 Segment
X4195 N4195 N4196 Segment
X4196 N4196 N4197 Segment
X4197 N4197 N4198 Segment
X4198 N4198 N4199 Segment
X4199 N4199 N4200 Segment
X4200 N4200 N4201 Segment
X4201 N4201 N4202 Segment
X4202 N4202 N4203 Segment
X4203 N4203 N4204 Segment
X4204 N4204 N4205 Segment
X4205 N4205 N4206 Segment
X4206 N4206 N4207 Segment
X4207 N4207 N4208 Segment
X4208 N4208 N4209 Segment
X4209 N4209 N4210 Segment
X4210 N4210 N4211 Segment
X4211 N4211 N4212 Segment
X4212 N4212 N4213 Segment
X4213 N4213 N4214 Segment
X4214 N4214 N4215 Segment
X4215 N4215 N4216 Segment
X4216 N4216 N4217 Segment
X4217 N4217 N4218 Segment
X4218 N4218 N4219 Segment
X4219 N4219 N4220 Segment
X4220 N4220 N4221 Segment
X4221 N4221 N4222 Segment
X4222 N4222 N4223 Segment
X4223 N4223 N4224 Segment
X4224 N4224 N4225 Segment
X4225 N4225 N4226 Segment
X4226 N4226 N4227 Segment
X4227 N4227 N4228 Segment
X4228 N4228 N4229 Segment
X4229 N4229 N4230 Segment
X4230 N4230 N4231 Segment
X4231 N4231 N4232 Segment
X4232 N4232 N4233 Segment
X4233 N4233 N4234 Segment
X4234 N4234 N4235 Segment
X4235 N4235 N4236 Segment
X4236 N4236 N4237 Segment
X4237 N4237 N4238 Segment
X4238 N4238 N4239 Segment
X4239 N4239 N4240 Segment
X4240 N4240 N4241 Segment
X4241 N4241 N4242 Segment
X4242 N4242 N4243 Segment
X4243 N4243 N4244 Segment
X4244 N4244 N4245 Segment
X4245 N4245 N4246 Segment
X4246 N4246 N4247 Segment
X4247 N4247 N4248 Segment
X4248 N4248 N4249 Segment
X4249 N4249 N4250 Segment
X4250 N4250 N4251 Segment
X4251 N4251 N4252 Segment
X4252 N4252 N4253 Segment
X4253 N4253 N4254 Segment
X4254 N4254 N4255 Segment
X4255 N4255 N4256 Segment
X4256 N4256 N4257 Segment
X4257 N4257 N4258 Segment
X4258 N4258 N4259 Segment
X4259 N4259 N4260 Segment
X4260 N4260 N4261 Segment
X4261 N4261 N4262 Segment
X4262 N4262 N4263 Segment
X4263 N4263 N4264 Segment
X4264 N4264 N4265 Segment
X4265 N4265 N4266 Segment
X4266 N4266 N4267 Segment
X4267 N4267 N4268 Segment
X4268 N4268 N4269 Segment
X4269 N4269 N4270 Segment
X4270 N4270 N4271 Segment
X4271 N4271 N4272 Segment
X4272 N4272 N4273 Segment
X4273 N4273 N4274 Segment
X4274 N4274 N4275 Segment
X4275 N4275 N4276 Segment
X4276 N4276 N4277 Segment
X4277 N4277 N4278 Segment
X4278 N4278 N4279 Segment
X4279 N4279 N4280 Segment
X4280 N4280 N4281 Segment
X4281 N4281 N4282 Segment
X4282 N4282 N4283 Segment
X4283 N4283 N4284 Segment
X4284 N4284 N4285 Segment
X4285 N4285 N4286 Segment
X4286 N4286 N4287 Segment
X4287 N4287 N4288 Segment
X4288 N4288 N4289 Segment
X4289 N4289 N4290 Segment
X4290 N4290 N4291 Segment
X4291 N4291 N4292 Segment
X4292 N4292 N4293 Segment
X4293 N4293 N4294 Segment
X4294 N4294 N4295 Segment
X4295 N4295 N4296 Segment
X4296 N4296 N4297 Segment
X4297 N4297 N4298 Segment
X4298 N4298 N4299 Segment
X4299 N4299 N4300 Segment
X4300 N4300 N4301 Segment
X4301 N4301 N4302 Segment
X4302 N4302 N4303 Segment
X4303 N4303 N4304 Segment
X4304 N4304 N4305 Segment
X4305 N4305 N4306 Segment
X4306 N4306 N4307 Segment
X4307 N4307 N4308 Segment
X4308 N4308 N4309 Segment
X4309 N4309 N4310 Segment
X4310 N4310 N4311 Segment
X4311 N4311 N4312 Segment
X4312 N4312 N4313 Segment
X4313 N4313 N4314 Segment
X4314 N4314 N4315 Segment
X4315 N4315 N4316 Segment
X4316 N4316 N4317 Segment
X4317 N4317 N4318 Segment
X4318 N4318 N4319 Segment
X4319 N4319 N4320 Segment
X4320 N4320 N4321 Segment
X4321 N4321 N4322 Segment
X4322 N4322 N4323 Segment
X4323 N4323 N4324 Segment
X4324 N4324 N4325 Segment
X4325 N4325 N4326 Segment
X4326 N4326 N4327 Segment
X4327 N4327 N4328 Segment
X4328 N4328 N4329 Segment
X4329 N4329 N4330 Segment
X4330 N4330 N4331 Segment
X4331 N4331 N4332 Segment
X4332 N4332 N4333 Segment
X4333 N4333 N4334 Segment
X4334 N4334 N4335 Segment
X4335 N4335 N4336 Segment
X4336 N4336 N4337 Segment
X4337 N4337 N4338 Segment
X4338 N4338 N4339 Segment
X4339 N4339 N4340 Segment
X4340 N4340 N4341 Segment
X4341 N4341 N4342 Segment
X4342 N4342 N4343 Segment
X4343 N4343 N4344 Segment
X4344 N4344 N4345 Segment
X4345 N4345 N4346 Segment
X4346 N4346 N4347 Segment
X4347 N4347 N4348 Segment
X4348 N4348 N4349 Segment
X4349 N4349 N4350 Segment
X4350 N4350 N4351 Segment
X4351 N4351 N4352 Segment
X4352 N4352 N4353 Segment
X4353 N4353 N4354 Segment
X4354 N4354 N4355 Segment
X4355 N4355 N4356 Segment
X4356 N4356 N4357 Segment
X4357 N4357 N4358 Segment
X4358 N4358 N4359 Segment
X4359 N4359 N4360 Segment
X4360 N4360 N4361 Segment
X4361 N4361 N4362 Segment
X4362 N4362 N4363 Segment
X4363 N4363 N4364 Segment
X4364 N4364 N4365 Segment
X4365 N4365 N4366 Segment
X4366 N4366 N4367 Segment
X4367 N4367 N4368 Segment
X4368 N4368 N4369 Segment
X4369 N4369 N4370 Segment
X4370 N4370 N4371 Segment
X4371 N4371 N4372 Segment
X4372 N4372 N4373 Segment
X4373 N4373 N4374 Segment
X4374 N4374 N4375 Segment
X4375 N4375 N4376 Segment
X4376 N4376 N4377 Segment
X4377 N4377 N4378 Segment
X4378 N4378 N4379 Segment
X4379 N4379 N4380 Segment
X4380 N4380 N4381 Segment
X4381 N4381 N4382 Segment
X4382 N4382 N4383 Segment
X4383 N4383 N4384 Segment
X4384 N4384 N4385 Segment
X4385 N4385 N4386 Segment
X4386 N4386 N4387 Segment
X4387 N4387 N4388 Segment
X4388 N4388 N4389 Segment
X4389 N4389 N4390 Segment
X4390 N4390 N4391 Segment
X4391 N4391 N4392 Segment
X4392 N4392 N4393 Segment
X4393 N4393 N4394 Segment
X4394 N4394 N4395 Segment
X4395 N4395 N4396 Segment
X4396 N4396 N4397 Segment
X4397 N4397 N4398 Segment
X4398 N4398 N4399 Segment
X4399 N4399 N4400 Segment
X4400 N4400 N4401 Segment
X4401 N4401 N4402 Segment
X4402 N4402 N4403 Segment
X4403 N4403 N4404 Segment
X4404 N4404 N4405 Segment
X4405 N4405 N4406 Segment
X4406 N4406 N4407 Segment
X4407 N4407 N4408 Segment
X4408 N4408 N4409 Segment
X4409 N4409 N4410 Segment
X4410 N4410 N4411 Segment
X4411 N4411 N4412 Segment
X4412 N4412 N4413 Segment
X4413 N4413 N4414 Segment
X4414 N4414 N4415 Segment
X4415 N4415 N4416 Segment
X4416 N4416 N4417 Segment
X4417 N4417 N4418 Segment
X4418 N4418 N4419 Segment
X4419 N4419 N4420 Segment
X4420 N4420 N4421 Segment
X4421 N4421 N4422 Segment
X4422 N4422 N4423 Segment
X4423 N4423 N4424 Segment
X4424 N4424 N4425 Segment
X4425 N4425 N4426 Segment
X4426 N4426 N4427 Segment
X4427 N4427 N4428 Segment
X4428 N4428 N4429 Segment
X4429 N4429 N4430 Segment
X4430 N4430 N4431 Segment
X4431 N4431 N4432 Segment
X4432 N4432 N4433 Segment
X4433 N4433 N4434 Segment
X4434 N4434 N4435 Segment
X4435 N4435 N4436 Segment
X4436 N4436 N4437 Segment
X4437 N4437 N4438 Segment
X4438 N4438 N4439 Segment
X4439 N4439 N4440 Segment
X4440 N4440 N4441 Segment
X4441 N4441 N4442 Segment
X4442 N4442 N4443 Segment
X4443 N4443 N4444 Segment
X4444 N4444 N4445 Segment
X4445 N4445 N4446 Segment
X4446 N4446 N4447 Segment
X4447 N4447 N4448 Segment
X4448 N4448 N4449 Segment
X4449 N4449 N4450 Segment
X4450 N4450 N4451 Segment
X4451 N4451 N4452 Segment
X4452 N4452 N4453 Segment
X4453 N4453 N4454 Segment
X4454 N4454 N4455 Segment
X4455 N4455 N4456 Segment
X4456 N4456 N4457 Segment
X4457 N4457 N4458 Segment
X4458 N4458 N4459 Segment
X4459 N4459 N4460 Segment
X4460 N4460 N4461 Segment
X4461 N4461 N4462 Segment
X4462 N4462 N4463 Segment
X4463 N4463 N4464 Segment
X4464 N4464 N4465 Segment
X4465 N4465 N4466 Segment
X4466 N4466 N4467 Segment
X4467 N4467 N4468 Segment
X4468 N4468 N4469 Segment
X4469 N4469 N4470 Segment
X4470 N4470 N4471 Segment
X4471 N4471 N4472 Segment
X4472 N4472 N4473 Segment
X4473 N4473 N4474 Segment
X4474 N4474 N4475 Segment
X4475 N4475 N4476 Segment
X4476 N4476 N4477 Segment
X4477 N4477 N4478 Segment
X4478 N4478 N4479 Segment
X4479 N4479 N4480 Segment
X4480 N4480 N4481 Segment
X4481 N4481 N4482 Segment
X4482 N4482 N4483 Segment
X4483 N4483 N4484 Segment
X4484 N4484 N4485 Segment
X4485 N4485 N4486 Segment
X4486 N4486 N4487 Segment
X4487 N4487 N4488 Segment
X4488 N4488 N4489 Segment
X4489 N4489 N4490 Segment
X4490 N4490 N4491 Segment
X4491 N4491 N4492 Segment
X4492 N4492 N4493 Segment
X4493 N4493 N4494 Segment
X4494 N4494 N4495 Segment
X4495 N4495 N4496 Segment
X4496 N4496 N4497 Segment
X4497 N4497 N4498 Segment
X4498 N4498 N4499 Segment
X4499 N4499 N4500 Segment
X4500 N4500 N4501 Segment
X4501 N4501 N4502 Segment
X4502 N4502 N4503 Segment
X4503 N4503 N4504 Segment
X4504 N4504 N4505 Segment
X4505 N4505 N4506 Segment
X4506 N4506 N4507 Segment
X4507 N4507 N4508 Segment
X4508 N4508 N4509 Segment
X4509 N4509 N4510 Segment
X4510 N4510 N4511 Segment
X4511 N4511 N4512 Segment
X4512 N4512 N4513 Segment
X4513 N4513 N4514 Segment
X4514 N4514 N4515 Segment
X4515 N4515 N4516 Segment
X4516 N4516 N4517 Segment
X4517 N4517 N4518 Segment
X4518 N4518 N4519 Segment
X4519 N4519 N4520 Segment
X4520 N4520 N4521 Segment
X4521 N4521 N4522 Segment
X4522 N4522 N4523 Segment
X4523 N4523 N4524 Segment
X4524 N4524 N4525 Segment
X4525 N4525 N4526 Segment
X4526 N4526 N4527 Segment
X4527 N4527 N4528 Segment
X4528 N4528 N4529 Segment
X4529 N4529 N4530 Segment
X4530 N4530 N4531 Segment
X4531 N4531 N4532 Segment
X4532 N4532 N4533 Segment
X4533 N4533 N4534 Segment
X4534 N4534 N4535 Segment
X4535 N4535 N4536 Segment
X4536 N4536 N4537 Segment
X4537 N4537 N4538 Segment
X4538 N4538 N4539 Segment
X4539 N4539 N4540 Segment
X4540 N4540 N4541 Segment
X4541 N4541 N4542 Segment
X4542 N4542 N4543 Segment
X4543 N4543 N4544 Segment
X4544 N4544 N4545 Segment
X4545 N4545 N4546 Segment
X4546 N4546 N4547 Segment
X4547 N4547 N4548 Segment
X4548 N4548 N4549 Segment
X4549 N4549 N4550 Segment
X4550 N4550 N4551 Segment
X4551 N4551 N4552 Segment
X4552 N4552 N4553 Segment
X4553 N4553 N4554 Segment
X4554 N4554 N4555 Segment
X4555 N4555 N4556 Segment
X4556 N4556 N4557 Segment
X4557 N4557 N4558 Segment
X4558 N4558 N4559 Segment
X4559 N4559 N4560 Segment
X4560 N4560 N4561 Segment
X4561 N4561 N4562 Segment
X4562 N4562 N4563 Segment
X4563 N4563 N4564 Segment
X4564 N4564 N4565 Segment
X4565 N4565 N4566 Segment
X4566 N4566 N4567 Segment
X4567 N4567 N4568 Segment
X4568 N4568 N4569 Segment
X4569 N4569 N4570 Segment
X4570 N4570 N4571 Segment
X4571 N4571 N4572 Segment
X4572 N4572 N4573 Segment
X4573 N4573 N4574 Segment
X4574 N4574 N4575 Segment
X4575 N4575 N4576 Segment
X4576 N4576 N4577 Segment
X4577 N4577 N4578 Segment
X4578 N4578 N4579 Segment
X4579 N4579 N4580 Segment
X4580 N4580 N4581 Segment
X4581 N4581 N4582 Segment
X4582 N4582 N4583 Segment
X4583 N4583 N4584 Segment
X4584 N4584 N4585 Segment
X4585 N4585 N4586 Segment
X4586 N4586 N4587 Segment
X4587 N4587 N4588 Segment
X4588 N4588 N4589 Segment
X4589 N4589 N4590 Segment
X4590 N4590 N4591 Segment
X4591 N4591 N4592 Segment
X4592 N4592 N4593 Segment
X4593 N4593 N4594 Segment
X4594 N4594 N4595 Segment
X4595 N4595 N4596 Segment
X4596 N4596 N4597 Segment
X4597 N4597 N4598 Segment
X4598 N4598 N4599 Segment
X4599 N4599 N4600 Segment
X4600 N4600 N4601 Segment
X4601 N4601 N4602 Segment
X4602 N4602 N4603 Segment
X4603 N4603 N4604 Segment
X4604 N4604 N4605 Segment
X4605 N4605 N4606 Segment
X4606 N4606 N4607 Segment
X4607 N4607 N4608 Segment
X4608 N4608 N4609 Segment
X4609 N4609 N4610 Segment
X4610 N4610 N4611 Segment
X4611 N4611 N4612 Segment
X4612 N4612 N4613 Segment
X4613 N4613 N4614 Segment
X4614 N4614 N4615 Segment
X4615 N4615 N4616 Segment
X4616 N4616 N4617 Segment
X4617 N4617 N4618 Segment
X4618 N4618 N4619 Segment
X4619 N4619 N4620 Segment
X4620 N4620 N4621 Segment
X4621 N4621 N4622 Segment
X4622 N4622 N4623 Segment
X4623 N4623 N4624 Segment
X4624 N4624 N4625 Segment
X4625 N4625 N4626 Segment
X4626 N4626 N4627 Segment
X4627 N4627 N4628 Segment
X4628 N4628 N4629 Segment
X4629 N4629 N4630 Segment
X4630 N4630 N4631 Segment
X4631 N4631 N4632 Segment
X4632 N4632 N4633 Segment
X4633 N4633 N4634 Segment
X4634 N4634 N4635 Segment
X4635 N4635 N4636 Segment
X4636 N4636 N4637 Segment
X4637 N4637 N4638 Segment
X4638 N4638 N4639 Segment
X4639 N4639 N4640 Segment
X4640 N4640 N4641 Segment
X4641 N4641 N4642 Segment
X4642 N4642 N4643 Segment
X4643 N4643 N4644 Segment
X4644 N4644 N4645 Segment
X4645 N4645 N4646 Segment
X4646 N4646 N4647 Segment
X4647 N4647 N4648 Segment
X4648 N4648 N4649 Segment
X4649 N4649 N4650 Segment
X4650 N4650 N4651 Segment
X4651 N4651 N4652 Segment
X4652 N4652 N4653 Segment
X4653 N4653 N4654 Segment
X4654 N4654 N4655 Segment
X4655 N4655 N4656 Segment
X4656 N4656 N4657 Segment
X4657 N4657 N4658 Segment
X4658 N4658 N4659 Segment
X4659 N4659 N4660 Segment
X4660 N4660 N4661 Segment
X4661 N4661 N4662 Segment
X4662 N4662 N4663 Segment
X4663 N4663 N4664 Segment
X4664 N4664 N4665 Segment
X4665 N4665 N4666 Segment
X4666 N4666 N4667 Segment
X4667 N4667 N4668 Segment
X4668 N4668 N4669 Segment
X4669 N4669 N4670 Segment
X4670 N4670 N4671 Segment
X4671 N4671 N4672 Segment
X4672 N4672 N4673 Segment
X4673 N4673 N4674 Segment
X4674 N4674 N4675 Segment
X4675 N4675 N4676 Segment
X4676 N4676 N4677 Segment
X4677 N4677 N4678 Segment
X4678 N4678 N4679 Segment
X4679 N4679 N4680 Segment
X4680 N4680 N4681 Segment
X4681 N4681 N4682 Segment
X4682 N4682 N4683 Segment
X4683 N4683 N4684 Segment
X4684 N4684 N4685 Segment
X4685 N4685 N4686 Segment
X4686 N4686 N4687 Segment
X4687 N4687 N4688 Segment
X4688 N4688 N4689 Segment
X4689 N4689 N4690 Segment
X4690 N4690 N4691 Segment
X4691 N4691 N4692 Segment
X4692 N4692 N4693 Segment
X4693 N4693 N4694 Segment
X4694 N4694 N4695 Segment
X4695 N4695 N4696 Segment
X4696 N4696 N4697 Segment
X4697 N4697 N4698 Segment
X4698 N4698 N4699 Segment
X4699 N4699 N4700 Segment
X4700 N4700 N4701 Segment
X4701 N4701 N4702 Segment
X4702 N4702 N4703 Segment
X4703 N4703 N4704 Segment
X4704 N4704 N4705 Segment
X4705 N4705 N4706 Segment
X4706 N4706 N4707 Segment
X4707 N4707 N4708 Segment
X4708 N4708 N4709 Segment
X4709 N4709 N4710 Segment
X4710 N4710 N4711 Segment
X4711 N4711 N4712 Segment
X4712 N4712 N4713 Segment
X4713 N4713 N4714 Segment
X4714 N4714 N4715 Segment
X4715 N4715 N4716 Segment
X4716 N4716 N4717 Segment
X4717 N4717 N4718 Segment
X4718 N4718 N4719 Segment
X4719 N4719 N4720 Segment
X4720 N4720 N4721 Segment
X4721 N4721 N4722 Segment
X4722 N4722 N4723 Segment
X4723 N4723 N4724 Segment
X4724 N4724 N4725 Segment
X4725 N4725 N4726 Segment
X4726 N4726 N4727 Segment
X4727 N4727 N4728 Segment
X4728 N4728 N4729 Segment
X4729 N4729 N4730 Segment
X4730 N4730 N4731 Segment
X4731 N4731 N4732 Segment
X4732 N4732 N4733 Segment
X4733 N4733 N4734 Segment
X4734 N4734 N4735 Segment
X4735 N4735 N4736 Segment
X4736 N4736 N4737 Segment
X4737 N4737 N4738 Segment
X4738 N4738 N4739 Segment
X4739 N4739 N4740 Segment
X4740 N4740 N4741 Segment
X4741 N4741 N4742 Segment
X4742 N4742 N4743 Segment
X4743 N4743 N4744 Segment
X4744 N4744 N4745 Segment
X4745 N4745 N4746 Segment
X4746 N4746 N4747 Segment
X4747 N4747 N4748 Segment
X4748 N4748 N4749 Segment
X4749 N4749 N4750 Segment
X4750 N4750 N4751 Segment
X4751 N4751 N4752 Segment
X4752 N4752 N4753 Segment
X4753 N4753 N4754 Segment
X4754 N4754 N4755 Segment
X4755 N4755 N4756 Segment
X4756 N4756 N4757 Segment
X4757 N4757 N4758 Segment
X4758 N4758 N4759 Segment
X4759 N4759 N4760 Segment
X4760 N4760 N4761 Segment
X4761 N4761 N4762 Segment
X4762 N4762 N4763 Segment
X4763 N4763 N4764 Segment
X4764 N4764 N4765 Segment
X4765 N4765 N4766 Segment
X4766 N4766 N4767 Segment
X4767 N4767 N4768 Segment
X4768 N4768 N4769 Segment
X4769 N4769 N4770 Segment
X4770 N4770 N4771 Segment
X4771 N4771 N4772 Segment
X4772 N4772 N4773 Segment
X4773 N4773 N4774 Segment
X4774 N4774 N4775 Segment
X4775 N4775 N4776 Segment
X4776 N4776 N4777 Segment
X4777 N4777 N4778 Segment
X4778 N4778 N4779 Segment
X4779 N4779 N4780 Segment
X4780 N4780 N4781 Segment
X4781 N4781 N4782 Segment
X4782 N4782 N4783 Segment
X4783 N4783 N4784 Segment
X4784 N4784 N4785 Segment
X4785 N4785 N4786 Segment
X4786 N4786 N4787 Segment
X4787 N4787 N4788 Segment
X4788 N4788 N4789 Segment
X4789 N4789 N4790 Segment
X4790 N4790 N4791 Segment
X4791 N4791 N4792 Segment
X4792 N4792 N4793 Segment
X4793 N4793 N4794 Segment
X4794 N4794 N4795 Segment
X4795 N4795 N4796 Segment
X4796 N4796 N4797 Segment
X4797 N4797 N4798 Segment
X4798 N4798 N4799 Segment
X4799 N4799 N4800 Segment
X4800 N4800 N4801 Segment
X4801 N4801 N4802 Segment
X4802 N4802 N4803 Segment
X4803 N4803 N4804 Segment
X4804 N4804 N4805 Segment
X4805 N4805 N4806 Segment
X4806 N4806 N4807 Segment
X4807 N4807 N4808 Segment
X4808 N4808 N4809 Segment
X4809 N4809 N4810 Segment
X4810 N4810 N4811 Segment
X4811 N4811 N4812 Segment
X4812 N4812 N4813 Segment
X4813 N4813 N4814 Segment
X4814 N4814 N4815 Segment
X4815 N4815 N4816 Segment
X4816 N4816 N4817 Segment
X4817 N4817 N4818 Segment
X4818 N4818 N4819 Segment
X4819 N4819 N4820 Segment
X4820 N4820 N4821 Segment
X4821 N4821 N4822 Segment
X4822 N4822 N4823 Segment
X4823 N4823 N4824 Segment
X4824 N4824 N4825 Segment
X4825 N4825 N4826 Segment
X4826 N4826 N4827 Segment
X4827 N4827 N4828 Segment
X4828 N4828 N4829 Segment
X4829 N4829 N4830 Segment
X4830 N4830 N4831 Segment
X4831 N4831 N4832 Segment
X4832 N4832 N4833 Segment
X4833 N4833 N4834 Segment
X4834 N4834 N4835 Segment
X4835 N4835 N4836 Segment
X4836 N4836 N4837 Segment
X4837 N4837 N4838 Segment
X4838 N4838 N4839 Segment
X4839 N4839 N4840 Segment
X4840 N4840 N4841 Segment
X4841 N4841 N4842 Segment
X4842 N4842 N4843 Segment
X4843 N4843 N4844 Segment
X4844 N4844 N4845 Segment
X4845 N4845 N4846 Segment
X4846 N4846 N4847 Segment
X4847 N4847 N4848 Segment
X4848 N4848 N4849 Segment
X4849 N4849 N4850 Segment
X4850 N4850 N4851 Segment
X4851 N4851 N4852 Segment
X4852 N4852 N4853 Segment
X4853 N4853 N4854 Segment
X4854 N4854 N4855 Segment
X4855 N4855 N4856 Segment
X4856 N4856 N4857 Segment
X4857 N4857 N4858 Segment
X4858 N4858 N4859 Segment
X4859 N4859 N4860 Segment
X4860 N4860 N4861 Segment
X4861 N4861 N4862 Segment
X4862 N4862 N4863 Segment
X4863 N4863 N4864 Segment
X4864 N4864 N4865 Segment
X4865 N4865 N4866 Segment
X4866 N4866 N4867 Segment
X4867 N4867 N4868 Segment
X4868 N4868 N4869 Segment
X4869 N4869 N4870 Segment
X4870 N4870 N4871 Segment
X4871 N4871 N4872 Segment
X4872 N4872 N4873 Segment
X4873 N4873 N4874 Segment
X4874 N4874 N4875 Segment
X4875 N4875 N4876 Segment
X4876 N4876 N4877 Segment
X4877 N4877 N4878 Segment
X4878 N4878 N4879 Segment
X4879 N4879 N4880 Segment
X4880 N4880 N4881 Segment
X4881 N4881 N4882 Segment
X4882 N4882 N4883 Segment
X4883 N4883 N4884 Segment
X4884 N4884 N4885 Segment
X4885 N4885 N4886 Segment
X4886 N4886 N4887 Segment
X4887 N4887 N4888 Segment
X4888 N4888 N4889 Segment
X4889 N4889 N4890 Segment
X4890 N4890 N4891 Segment
X4891 N4891 N4892 Segment
X4892 N4892 N4893 Segment
X4893 N4893 N4894 Segment
X4894 N4894 N4895 Segment
X4895 N4895 N4896 Segment
X4896 N4896 N4897 Segment
X4897 N4897 N4898 Segment
X4898 N4898 N4899 Segment
X4899 N4899 N4900 Segment
X4900 N4900 N4901 Segment
X4901 N4901 N4902 Segment
X4902 N4902 N4903 Segment
X4903 N4903 N4904 Segment
X4904 N4904 N4905 Segment
X4905 N4905 N4906 Segment
X4906 N4906 N4907 Segment
X4907 N4907 N4908 Segment
X4908 N4908 N4909 Segment
X4909 N4909 N4910 Segment
X4910 N4910 N4911 Segment
X4911 N4911 N4912 Segment
X4912 N4912 N4913 Segment
X4913 N4913 N4914 Segment
X4914 N4914 N4915 Segment
X4915 N4915 N4916 Segment
X4916 N4916 N4917 Segment
X4917 N4917 N4918 Segment
X4918 N4918 N4919 Segment
X4919 N4919 N4920 Segment
X4920 N4920 N4921 Segment
X4921 N4921 N4922 Segment
X4922 N4922 N4923 Segment
X4923 N4923 N4924 Segment
X4924 N4924 N4925 Segment
X4925 N4925 N4926 Segment
X4926 N4926 N4927 Segment
X4927 N4927 N4928 Segment
X4928 N4928 N4929 Segment
X4929 N4929 N4930 Segment
X4930 N4930 N4931 Segment
X4931 N4931 N4932 Segment
X4932 N4932 N4933 Segment
X4933 N4933 N4934 Segment
X4934 N4934 N4935 Segment
X4935 N4935 N4936 Segment
X4936 N4936 N4937 Segment
X4937 N4937 N4938 Segment
X4938 N4938 N4939 Segment
X4939 N4939 N4940 Segment
X4940 N4940 N4941 Segment
X4941 N4941 N4942 Segment
X4942 N4942 N4943 Segment
X4943 N4943 N4944 Segment
X4944 N4944 N4945 Segment
X4945 N4945 N4946 Segment
X4946 N4946 N4947 Segment
X4947 N4947 N4948 Segment
X4948 N4948 N4949 Segment
X4949 N4949 N4950 Segment
X4950 N4950 N4951 Segment
X4951 N4951 N4952 Segment
X4952 N4952 N4953 Segment
X4953 N4953 N4954 Segment
X4954 N4954 N4955 Segment
X4955 N4955 N4956 Segment
X4956 N4956 N4957 Segment
X4957 N4957 N4958 Segment
X4958 N4958 N4959 Segment
X4959 N4959 N4960 Segment
X4960 N4960 N4961 Segment
X4961 N4961 N4962 Segment
X4962 N4962 N4963 Segment
X4963 N4963 N4964 Segment
X4964 N4964 N4965 Segment
X4965 N4965 N4966 Segment
X4966 N4966 N4967 Segment
X4967 N4967 N4968 Segment
X4968 N4968 N4969 Segment
X4969 N4969 N4970 Segment
X4970 N4970 N4971 Segment
X4971 N4971 N4972 Segment
X4972 N4972 N4973 Segment
X4973 N4973 N4974 Segment
X4974 N4974 N4975 Segment
X4975 N4975 N4976 Segment
X4976 N4976 N4977 Segment
X4977 N4977 N4978 Segment
X4978 N4978 N4979 Segment
X4979 N4979 N4980 Segment
X4980 N4980 N4981 Segment
X4981 N4981 N4982 Segment
X4982 N4982 N4983 Segment
X4983 N4983 N4984 Segment
X4984 N4984 N4985 Segment
X4985 N4985 N4986 Segment
X4986 N4986 N4987 Segment
X4987 N4987 N4988 Segment
X4988 N4988 N4989 Segment
X4989 N4989 N4990 Segment
X4990 N4990 N4991 Segment
X4991 N4991 N4992 Segment
X4992 N4992 N4993 Segment
X4993 N4993 N4994 Segment
X4994 N4994 N4995 Segment
X4995 N4995 N4996 Segment
X4996 N4996 N4997 Segment
X4997 N4997 N4998 Segment
X4998 N4998 N4999 Segment
X4999 N4999 N5000 Segment
X5000 N5000 N5001 Segment
X5001 N5001 N5002 Segment
X5002 N5002 N5003 Segment
X5003 N5003 N5004 Segment
X5004 N5004 N5005 Segment
X5005 N5005 N5006 Segment
X5006 N5006 N5007 Segment
X5007 N5007 N5008 Segment
X5008 N5008 N5009 Segment
X5009 N5009 N5010 Segment
X5010 N5010 N5011 Segment
X5011 N5011 N5012 Segment
X5012 N5012 N5013 Segment
X5013 N5013 N5014 Segment
X5014 N5014 N5015 Segment
X5015 N5015 N5016 Segment
X5016 N5016 N5017 Segment
X5017 N5017 N5018 Segment
X5018 N5018 N5019 Segment
X5019 N5019 N5020 Segment
X5020 N5020 N5021 Segment
X5021 N5021 N5022 Segment
X5022 N5022 N5023 Segment
X5023 N5023 N5024 Segment
X5024 N5024 N5025 Segment
X5025 N5025 N5026 Segment
X5026 N5026 N5027 Segment
X5027 N5027 N5028 Segment
X5028 N5028 N5029 Segment
X5029 N5029 N5030 Segment
X5030 N5030 N5031 Segment
X5031 N5031 N5032 Segment
X5032 N5032 N5033 Segment
X5033 N5033 N5034 Segment
X5034 N5034 N5035 Segment
X5035 N5035 N5036 Segment
X5036 N5036 N5037 Segment
X5037 N5037 N5038 Segment
X5038 N5038 N5039 Segment
X5039 N5039 N5040 Segment
X5040 N5040 N5041 Segment
X5041 N5041 N5042 Segment
X5042 N5042 N5043 Segment
X5043 N5043 N5044 Segment
X5044 N5044 N5045 Segment
X5045 N5045 N5046 Segment
X5046 N5046 N5047 Segment
X5047 N5047 N5048 Segment
X5048 N5048 N5049 Segment
X5049 N5049 N5050 Segment
X5050 N5050 N5051 Segment
X5051 N5051 N5052 Segment
X5052 N5052 N5053 Segment
X5053 N5053 N5054 Segment
X5054 N5054 N5055 Segment
X5055 N5055 N5056 Segment
X5056 N5056 N5057 Segment
X5057 N5057 N5058 Segment
X5058 N5058 N5059 Segment
X5059 N5059 N5060 Segment
X5060 N5060 N5061 Segment
X5061 N5061 N5062 Segment
X5062 N5062 N5063 Segment
X5063 N5063 N5064 Segment
X5064 N5064 N5065 Segment
X5065 N5065 N5066 Segment
X5066 N5066 N5067 Segment
X5067 N5067 N5068 Segment
X5068 N5068 N5069 Segment
X5069 N5069 N5070 Segment
X5070 N5070 N5071 Segment
X5071 N5071 N5072 Segment
X5072 N5072 N5073 Segment
X5073 N5073 N5074 Segment
X5074 N5074 N5075 Segment
X5075 N5075 N5076 Segment
X5076 N5076 N5077 Segment
X5077 N5077 N5078 Segment
X5078 N5078 N5079 Segment
X5079 N5079 N5080 Segment
X5080 N5080 N5081 Segment
X5081 N5081 N5082 Segment
X5082 N5082 N5083 Segment
X5083 N5083 N5084 Segment
X5084 N5084 N5085 Segment
X5085 N5085 N5086 Segment
X5086 N5086 N5087 Segment
X5087 N5087 N5088 Segment
X5088 N5088 N5089 Segment
X5089 N5089 N5090 Segment
X5090 N5090 N5091 Segment
X5091 N5091 N5092 Segment
X5092 N5092 N5093 Segment
X5093 N5093 N5094 Segment
X5094 N5094 N5095 Segment
X5095 N5095 N5096 Segment
X5096 N5096 N5097 Segment
X5097 N5097 N5098 Segment
X5098 N5098 N5099 Segment
X5099 N5099 N5100 Segment
X5100 N5100 N5101 Segment
X5101 N5101 N5102 Segment
X5102 N5102 N5103 Segment
X5103 N5103 N5104 Segment
X5104 N5104 N5105 Segment
X5105 N5105 N5106 Segment
X5106 N5106 N5107 Segment
X5107 N5107 N5108 Segment
X5108 N5108 N5109 Segment
X5109 N5109 N5110 Segment
X5110 N5110 N5111 Segment
X5111 N5111 N5112 Segment
X5112 N5112 N5113 Segment
X5113 N5113 N5114 Segment
X5114 N5114 N5115 Segment
X5115 N5115 N5116 Segment
X5116 N5116 N5117 Segment
X5117 N5117 N5118 Segment
X5118 N5118 N5119 Segment
X5119 N5119 N5120 Segment
X5120 N5120 N5121 Segment
X5121 N5121 N5122 Segment
X5122 N5122 N5123 Segment
X5123 N5123 N5124 Segment
X5124 N5124 N5125 Segment
X5125 N5125 N5126 Segment
X5126 N5126 N5127 Segment
X5127 N5127 N5128 Segment
X5128 N5128 N5129 Segment
X5129 N5129 N5130 Segment
X5130 N5130 N5131 Segment
X5131 N5131 N5132 Segment
X5132 N5132 N5133 Segment
X5133 N5133 N5134 Segment
X5134 N5134 N5135 Segment
X5135 N5135 N5136 Segment
X5136 N5136 N5137 Segment
X5137 N5137 N5138 Segment
X5138 N5138 N5139 Segment
X5139 N5139 N5140 Segment
X5140 N5140 N5141 Segment
X5141 N5141 N5142 Segment
X5142 N5142 N5143 Segment
X5143 N5143 N5144 Segment
X5144 N5144 N5145 Segment
X5145 N5145 N5146 Segment
X5146 N5146 N5147 Segment
X5147 N5147 N5148 Segment
X5148 N5148 N5149 Segment
X5149 N5149 N5150 Segment
X5150 N5150 N5151 Segment
X5151 N5151 N5152 Segment
X5152 N5152 N5153 Segment
X5153 N5153 N5154 Segment
X5154 N5154 N5155 Segment
X5155 N5155 N5156 Segment
X5156 N5156 N5157 Segment
X5157 N5157 N5158 Segment
X5158 N5158 N5159 Segment
X5159 N5159 N5160 Segment
X5160 N5160 N5161 Segment
X5161 N5161 N5162 Segment
X5162 N5162 N5163 Segment
X5163 N5163 N5164 Segment
X5164 N5164 N5165 Segment
X5165 N5165 N5166 Segment
X5166 N5166 N5167 Segment
X5167 N5167 N5168 Segment
X5168 N5168 N5169 Segment
X5169 N5169 N5170 Segment
X5170 N5170 N5171 Segment
X5171 N5171 N5172 Segment
X5172 N5172 N5173 Segment
X5173 N5173 N5174 Segment
X5174 N5174 N5175 Segment
X5175 N5175 N5176 Segment
X5176 N5176 N5177 Segment
X5177 N5177 N5178 Segment
X5178 N5178 N5179 Segment
X5179 N5179 N5180 Segment
X5180 N5180 N5181 Segment
X5181 N5181 N5182 Segment
X5182 N5182 N5183 Segment
X5183 N5183 N5184 Segment
X5184 N5184 N5185 Segment
X5185 N5185 N5186 Segment
X5186 N5186 N5187 Segment
X5187 N5187 N5188 Segment
X5188 N5188 N5189 Segment
X5189 N5189 N5190 Segment
X5190 N5190 N5191 Segment
X5191 N5191 N5192 Segment
X5192 N5192 N5193 Segment
X5193 N5193 N5194 Segment
X5194 N5194 N5195 Segment
X5195 N5195 N5196 Segment
X5196 N5196 N5197 Segment
X5197 N5197 N5198 Segment
X5198 N5198 N5199 Segment
X5199 N5199 N5200 Segment
X5200 N5200 N5201 Segment
X5201 N5201 N5202 Segment
X5202 N5202 N5203 Segment
X5203 N5203 N5204 Segment
X5204 N5204 N5205 Segment
X5205 N5205 N5206 Segment
X5206 N5206 N5207 Segment
X5207 N5207 N5208 Segment
X5208 N5208 N5209 Segment
X5209 N5209 N5210 Segment
X5210 N5210 N5211 Segment
X5211 N5211 N5212 Segment
X5212 N5212 N5213 Segment
X5213 N5213 N5214 Segment
X5214 N5214 N5215 Segment
X5215 N5215 N5216 Segment
X5216 N5216 N5217 Segment
X5217 N5217 N5218 Segment
X5218 N5218 N5219 Segment
X5219 N5219 N5220 Segment
X5220 N5220 N5221 Segment
X5221 N5221 N5222 Segment
X5222 N5222 N5223 Segment
X5223 N5223 N5224 Segment
X5224 N5224 N5225 Segment
X5225 N5225 N5226 Segment
X5226 N5226 N5227 Segment
X5227 N5227 N5228 Segment
X5228 N5228 N5229 Segment
X5229 N5229 N5230 Segment
X5230 N5230 N5231 Segment
X5231 N5231 N5232 Segment
X5232 N5232 N5233 Segment
X5233 N5233 N5234 Segment
X5234 N5234 N5235 Segment
X5235 N5235 N5236 Segment
X5236 N5236 N5237 Segment
X5237 N5237 N5238 Segment
X5238 N5238 N5239 Segment
X5239 N5239 N5240 Segment
X5240 N5240 N5241 Segment
X5241 N5241 N5242 Segment
X5242 N5242 N5243 Segment
X5243 N5243 N5244 Segment
X5244 N5244 N5245 Segment
X5245 N5245 N5246 Segment
X5246 N5246 N5247 Segment
X5247 N5247 N5248 Segment
X5248 N5248 N5249 Segment
X5249 N5249 N5250 Segment
X5250 N5250 N5251 Segment
X5251 N5251 N5252 Segment
X5252 N5252 N5253 Segment
X5253 N5253 N5254 Segment
X5254 N5254 N5255 Segment
X5255 N5255 N5256 Segment
X5256 N5256 N5257 Segment
X5257 N5257 N5258 Segment
X5258 N5258 N5259 Segment
X5259 N5259 N5260 Segment
X5260 N5260 N5261 Segment
X5261 N5261 N5262 Segment
X5262 N5262 N5263 Segment
X5263 N5263 N5264 Segment
X5264 N5264 N5265 Segment
X5265 N5265 N5266 Segment
X5266 N5266 N5267 Segment
X5267 N5267 N5268 Segment
X5268 N5268 N5269 Segment
X5269 N5269 N5270 Segment
X5270 N5270 N5271 Segment
X5271 N5271 N5272 Segment
X5272 N5272 N5273 Segment
X5273 N5273 N5274 Segment
X5274 N5274 N5275 Segment
X5275 N5275 N5276 Segment
X5276 N5276 N5277 Segment
X5277 N5277 N5278 Segment
X5278 N5278 N5279 Segment
X5279 N5279 N5280 Segment
X5280 N5280 N5281 Segment
X5281 N5281 N5282 Segment
X5282 N5282 N5283 Segment
X5283 N5283 N5284 Segment
X5284 N5284 N5285 Segment
X5285 N5285 N5286 Segment
X5286 N5286 N5287 Segment
X5287 N5287 N5288 Segment
X5288 N5288 N5289 Segment
X5289 N5289 N5290 Segment
X5290 N5290 N5291 Segment
X5291 N5291 N5292 Segment
X5292 N5292 N5293 Segment
X5293 N5293 N5294 Segment
X5294 N5294 N5295 Segment
X5295 N5295 N5296 Segment
X5296 N5296 N5297 Segment
X5297 N5297 N5298 Segment
X5298 N5298 N5299 Segment
X5299 N5299 N5300 Segment
X5300 N5300 N5301 Segment
X5301 N5301 N5302 Segment
X5302 N5302 N5303 Segment
X5303 N5303 N5304 Segment
X5304 N5304 N5305 Segment
X5305 N5305 N5306 Segment
X5306 N5306 N5307 Segment
X5307 N5307 N5308 Segment
X5308 N5308 N5309 Segment
X5309 N5309 N5310 Segment
X5310 N5310 N5311 Segment
X5311 N5311 N5312 Segment
X5312 N5312 N5313 Segment
X5313 N5313 N5314 Segment
X5314 N5314 N5315 Segment
X5315 N5315 N5316 Segment
X5316 N5316 N5317 Segment
X5317 N5317 N5318 Segment
X5318 N5318 N5319 Segment
X5319 N5319 N5320 Segment
X5320 N5320 N5321 Segment
X5321 N5321 N5322 Segment
X5322 N5322 N5323 Segment
X5323 N5323 N5324 Segment
X5324 N5324 N5325 Segment
X5325 N5325 N5326 Segment
X5326 N5326 N5327 Segment
X5327 N5327 N5328 Segment
X5328 N5328 N5329 Segment
X5329 N5329 N5330 Segment
X5330 N5330 N5331 Segment
X5331 N5331 N5332 Segment
X5332 N5332 N5333 Segment
X5333 N5333 N5334 Segment
X5334 N5334 N5335 Segment
X5335 N5335 N5336 Segment
X5336 N5336 N5337 Segment
X5337 N5337 N5338 Segment
X5338 N5338 N5339 Segment
X5339 N5339 N5340 Segment
X5340 N5340 N5341 Segment
X5341 N5341 N5342 Segment
X5342 N5342 N5343 Segment
X5343 N5343 N5344 Segment
X5344 N5344 N5345 Segment
X5345 N5345 N5346 Segment
X5346 N5346 N5347 Segment
X5347 N5347 N5348 Segment
X5348 N5348 N5349 Segment
X5349 N5349 N5350 Segment
X5350 N5350 N5351 Segment
X5351 N5351 N5352 Segment
X5352 N5352 N5353 Segment
X5353 N5353 N5354 Segment
X5354 N5354 N5355 Segment
X5355 N5355 N5356 Segment
X5356 N5356 N5357 Segment
X5357 N5357 N5358 Segment
X5358 N5358 N5359 Segment
X5359 N5359 N5360 Segment
X5360 N5360 N5361 Segment
X5361 N5361 N5362 Segment
X5362 N5362 N5363 Segment
X5363 N5363 N5364 Segment
X5364 N5364 N5365 Segment
X5365 N5365 N5366 Segment
X5366 N5366 N5367 Segment
X5367 N5367 N5368 Segment
X5368 N5368 N5369 Segment
X5369 N5369 N5370 Segment
X5370 N5370 N5371 Segment
X5371 N5371 N5372 Segment
X5372 N5372 N5373 Segment
X5373 N5373 N5374 Segment
X5374 N5374 N5375 Segment
X5375 N5375 N5376 Segment
X5376 N5376 N5377 Segment
X5377 N5377 N5378 Segment
X5378 N5378 N5379 Segment
X5379 N5379 N5380 Segment
X5380 N5380 N5381 Segment
X5381 N5381 N5382 Segment
X5382 N5382 N5383 Segment
X5383 N5383 N5384 Segment
X5384 N5384 N5385 Segment
X5385 N5385 N5386 Segment
X5386 N5386 N5387 Segment
X5387 N5387 N5388 Segment
X5388 N5388 N5389 Segment
X5389 N5389 N5390 Segment
X5390 N5390 N5391 Segment
X5391 N5391 N5392 Segment
X5392 N5392 N5393 Segment
X5393 N5393 N5394 Segment
X5394 N5394 N5395 Segment
X5395 N5395 N5396 Segment
X5396 N5396 N5397 Segment
X5397 N5397 N5398 Segment
X5398 N5398 N5399 Segment
X5399 N5399 N5400 Segment
X5400 N5400 N5401 Segment
X5401 N5401 N5402 Segment
X5402 N5402 N5403 Segment
X5403 N5403 N5404 Segment
X5404 N5404 N5405 Segment
X5405 N5405 N5406 Segment
X5406 N5406 N5407 Segment
X5407 N5407 N5408 Segment
X5408 N5408 N5409 Segment
X5409 N5409 N5410 Segment
X5410 N5410 N5411 Segment
X5411 N5411 N5412 Segment
X5412 N5412 N5413 Segment
X5413 N5413 N5414 Segment
X5414 N5414 N5415 Segment
X5415 N5415 N5416 Segment
X5416 N5416 N5417 Segment
X5417 N5417 N5418 Segment
X5418 N5418 N5419 Segment
X5419 N5419 N5420 Segment
X5420 N5420 N5421 Segment
X5421 N5421 N5422 Segment
X5422 N5422 N5423 Segment
X5423 N5423 N5424 Segment
X5424 N5424 N5425 Segment
X5425 N5425 N5426 Segment
X5426 N5426 N5427 Segment
X5427 N5427 N5428 Segment
X5428 N5428 N5429 Segment
X5429 N5429 N5430 Segment
X5430 N5430 N5431 Segment
X5431 N5431 N5432 Segment
X5432 N5432 N5433 Segment
X5433 N5433 N5434 Segment
X5434 N5434 N5435 Segment
X5435 N5435 N5436 Segment
X5436 N5436 N5437 Segment
X5437 N5437 N5438 Segment
X5438 N5438 N5439 Segment
X5439 N5439 N5440 Segment
X5440 N5440 N5441 Segment
X5441 N5441 N5442 Segment
X5442 N5442 N5443 Segment
X5443 N5443 N5444 Segment
X5444 N5444 N5445 Segment
X5445 N5445 N5446 Segment
X5446 N5446 N5447 Segment
X5447 N5447 N5448 Segment
X5448 N5448 N5449 Segment
X5449 N5449 N5450 Segment
X5450 N5450 N5451 Segment
X5451 N5451 N5452 Segment
X5452 N5452 N5453 Segment
X5453 N5453 N5454 Segment
X5454 N5454 N5455 Segment
X5455 N5455 N5456 Segment
X5456 N5456 N5457 Segment
X5457 N5457 N5458 Segment
X5458 N5458 N5459 Segment
X5459 N5459 N5460 Segment
X5460 N5460 N5461 Segment
X5461 N5461 N5462 Segment
X5462 N5462 N5463 Segment
X5463 N5463 N5464 Segment
X5464 N5464 N5465 Segment
X5465 N5465 N5466 Segment
X5466 N5466 N5467 Segment
X5467 N5467 N5468 Segment
X5468 N5468 N5469 Segment
X5469 N5469 N5470 Segment
X5470 N5470 N5471 Segment
X5471 N5471 N5472 Segment
X5472 N5472 N5473 Segment
X5473 N5473 N5474 Segment
X5474 N5474 N5475 Segment
X5475 N5475 N5476 Segment
X5476 N5476 N5477 Segment
X5477 N5477 N5478 Segment
X5478 N5478 N5479 Segment
X5479 N5479 N5480 Segment
X5480 N5480 N5481 Segment
X5481 N5481 N5482 Segment
X5482 N5482 N5483 Segment
X5483 N5483 N5484 Segment
X5484 N5484 N5485 Segment
X5485 N5485 N5486 Segment
X5486 N5486 N5487 Segment
X5487 N5487 N5488 Segment
X5488 N5488 N5489 Segment
X5489 N5489 N5490 Segment
X5490 N5490 N5491 Segment
X5491 N5491 N5492 Segment
X5492 N5492 N5493 Segment
X5493 N5493 N5494 Segment
X5494 N5494 N5495 Segment
X5495 N5495 N5496 Segment
X5496 N5496 N5497 Segment
X5497 N5497 N5498 Segment
X5498 N5498 N5499 Segment
X5499 N5499 N5500 Segment
X5500 N5500 N5501 Segment
X5501 N5501 N5502 Segment
X5502 N5502 N5503 Segment
X5503 N5503 N5504 Segment
X5504 N5504 N5505 Segment
X5505 N5505 N5506 Segment
X5506 N5506 N5507 Segment
X5507 N5507 N5508 Segment
X5508 N5508 N5509 Segment
X5509 N5509 N5510 Segment
X5510 N5510 N5511 Segment
X5511 N5511 N5512 Segment
X5512 N5512 N5513 Segment
X5513 N5513 N5514 Segment
X5514 N5514 N5515 Segment
X5515 N5515 N5516 Segment
X5516 N5516 N5517 Segment
X5517 N5517 N5518 Segment
X5518 N5518 N5519 Segment
X5519 N5519 N5520 Segment
X5520 N5520 N5521 Segment
X5521 N5521 N5522 Segment
X5522 N5522 N5523 Segment
X5523 N5523 N5524 Segment
X5524 N5524 N5525 Segment
X5525 N5525 N5526 Segment
X5526 N5526 N5527 Segment
X5527 N5527 N5528 Segment
X5528 N5528 N5529 Segment
X5529 N5529 N5530 Segment
X5530 N5530 N5531 Segment
X5531 N5531 N5532 Segment
X5532 N5532 N5533 Segment
X5533 N5533 N5534 Segment
X5534 N5534 N5535 Segment
X5535 N5535 N5536 Segment
X5536 N5536 N5537 Segment
X5537 N5537 N5538 Segment
X5538 N5538 N5539 Segment
X5539 N5539 N5540 Segment
X5540 N5540 N5541 Segment
X5541 N5541 N5542 Segment
X5542 N5542 N5543 Segment
X5543 N5543 N5544 Segment
X5544 N5544 N5545 Segment
X5545 N5545 N5546 Segment
X5546 N5546 N5547 Segment
X5547 N5547 N5548 Segment
X5548 N5548 N5549 Segment
X5549 N5549 N5550 Segment
X5550 N5550 N5551 Segment
X5551 N5551 N5552 Segment
X5552 N5552 N5553 Segment
X5553 N5553 N5554 Segment
X5554 N5554 N5555 Segment
X5555 N5555 N5556 Segment
X5556 N5556 N5557 Segment
X5557 N5557 N5558 Segment
X5558 N5558 N5559 Segment
X5559 N5559 N5560 Segment
X5560 N5560 N5561 Segment
X5561 N5561 N5562 Segment
X5562 N5562 N5563 Segment
X5563 N5563 N5564 Segment
X5564 N5564 N5565 Segment
X5565 N5565 N5566 Segment
X5566 N5566 N5567 Segment
X5567 N5567 N5568 Segment
X5568 N5568 N5569 Segment
X5569 N5569 N5570 Segment
X5570 N5570 N5571 Segment
X5571 N5571 N5572 Segment
X5572 N5572 N5573 Segment
X5573 N5573 N5574 Segment
X5574 N5574 N5575 Segment
X5575 N5575 N5576 Segment
X5576 N5576 N5577 Segment
X5577 N5577 N5578 Segment
X5578 N5578 N5579 Segment
X5579 N5579 N5580 Segment
X5580 N5580 N5581 Segment
X5581 N5581 N5582 Segment
X5582 N5582 N5583 Segment
X5583 N5583 N5584 Segment
X5584 N5584 N5585 Segment
X5585 N5585 N5586 Segment
X5586 N5586 N5587 Segment
X5587 N5587 N5588 Segment
X5588 N5588 N5589 Segment
X5589 N5589 N5590 Segment
X5590 N5590 N5591 Segment
X5591 N5591 N5592 Segment
X5592 N5592 N5593 Segment
X5593 N5593 N5594 Segment
X5594 N5594 N5595 Segment
X5595 N5595 N5596 Segment
X5596 N5596 N5597 Segment
X5597 N5597 N5598 Segment
X5598 N5598 N5599 Segment
X5599 N5599 N5600 Segment
X5600 N5600 N5601 Segment
X5601 N5601 N5602 Segment
X5602 N5602 N5603 Segment
X5603 N5603 N5604 Segment
X5604 N5604 N5605 Segment
X5605 N5605 N5606 Segment
X5606 N5606 N5607 Segment
X5607 N5607 N5608 Segment
X5608 N5608 N5609 Segment
X5609 N5609 N5610 Segment
X5610 N5610 N5611 Segment
X5611 N5611 N5612 Segment
X5612 N5612 N5613 Segment
X5613 N5613 N5614 Segment
X5614 N5614 N5615 Segment
X5615 N5615 N5616 Segment
X5616 N5616 N5617 Segment
X5617 N5617 N5618 Segment
X5618 N5618 N5619 Segment
X5619 N5619 N5620 Segment
X5620 N5620 N5621 Segment
X5621 N5621 N5622 Segment
X5622 N5622 N5623 Segment
X5623 N5623 N5624 Segment
X5624 N5624 N5625 Segment
X5625 N5625 N5626 Segment
X5626 N5626 N5627 Segment
X5627 N5627 N5628 Segment
X5628 N5628 N5629 Segment
X5629 N5629 N5630 Segment
X5630 N5630 N5631 Segment
X5631 N5631 N5632 Segment
X5632 N5632 N5633 Segment
X5633 N5633 N5634 Segment
X5634 N5634 N5635 Segment
X5635 N5635 N5636 Segment
X5636 N5636 N5637 Segment
X5637 N5637 N5638 Segment
X5638 N5638 N5639 Segment
X5639 N5639 N5640 Segment
X5640 N5640 N5641 Segment
X5641 N5641 N5642 Segment
X5642 N5642 N5643 Segment
X5643 N5643 N5644 Segment
X5644 N5644 N5645 Segment
X5645 N5645 N5646 Segment
X5646 N5646 N5647 Segment
X5647 N5647 N5648 Segment
X5648 N5648 N5649 Segment
X5649 N5649 N5650 Segment
X5650 N5650 N5651 Segment
X5651 N5651 N5652 Segment
X5652 N5652 N5653 Segment
X5653 N5653 N5654 Segment
X5654 N5654 N5655 Segment
X5655 N5655 N5656 Segment
X5656 N5656 N5657 Segment
X5657 N5657 N5658 Segment
X5658 N5658 N5659 Segment
X5659 N5659 N5660 Segment
X5660 N5660 N5661 Segment
X5661 N5661 N5662 Segment
X5662 N5662 N5663 Segment
X5663 N5663 N5664 Segment
X5664 N5664 N5665 Segment
X5665 N5665 N5666 Segment
X5666 N5666 N5667 Segment
X5667 N5667 N5668 Segment
X5668 N5668 N5669 Segment
X5669 N5669 N5670 Segment
X5670 N5670 N5671 Segment
X5671 N5671 N5672 Segment
X5672 N5672 N5673 Segment
X5673 N5673 N5674 Segment
X5674 N5674 N5675 Segment
X5675 N5675 N5676 Segment
X5676 N5676 N5677 Segment
X5677 N5677 N5678 Segment
X5678 N5678 N5679 Segment
X5679 N5679 N5680 Segment
X5680 N5680 N5681 Segment
X5681 N5681 N5682 Segment
X5682 N5682 N5683 Segment
X5683 N5683 N5684 Segment
X5684 N5684 N5685 Segment
X5685 N5685 N5686 Segment
X5686 N5686 N5687 Segment
X5687 N5687 N5688 Segment
X5688 N5688 N5689 Segment
X5689 N5689 N5690 Segment
X5690 N5690 N5691 Segment
X5691 N5691 N5692 Segment
X5692 N5692 N5693 Segment
X5693 N5693 N5694 Segment
X5694 N5694 N5695 Segment
X5695 N5695 N5696 Segment
X5696 N5696 N5697 Segment
X5697 N5697 N5698 Segment
X5698 N5698 N5699 Segment
X5699 N5699 N5700 Segment
X5700 N5700 N5701 Segment
X5701 N5701 N5702 Segment
X5702 N5702 N5703 Segment
X5703 N5703 N5704 Segment
X5704 N5704 N5705 Segment
X5705 N5705 N5706 Segment
X5706 N5706 N5707 Segment
X5707 N5707 N5708 Segment
X5708 N5708 N5709 Segment
X5709 N5709 N5710 Segment
X5710 N5710 N5711 Segment
X5711 N5711 N5712 Segment
X5712 N5712 N5713 Segment
X5713 N5713 N5714 Segment
X5714 N5714 N5715 Segment
X5715 N5715 N5716 Segment
X5716 N5716 N5717 Segment
X5717 N5717 N5718 Segment
X5718 N5718 N5719 Segment
X5719 N5719 N5720 Segment
X5720 N5720 N5721 Segment
X5721 N5721 N5722 Segment
X5722 N5722 N5723 Segment
X5723 N5723 N5724 Segment
X5724 N5724 N5725 Segment
X5725 N5725 N5726 Segment
X5726 N5726 N5727 Segment
X5727 N5727 N5728 Segment
X5728 N5728 N5729 Segment
X5729 N5729 N5730 Segment
X5730 N5730 N5731 Segment
X5731 N5731 N5732 Segment
X5732 N5732 N5733 Segment
X5733 N5733 N5734 Segment
X5734 N5734 N5735 Segment
X5735 N5735 N5736 Segment
X5736 N5736 N5737 Segment
X5737 N5737 N5738 Segment
X5738 N5738 N5739 Segment
X5739 N5739 N5740 Segment
X5740 N5740 N5741 Segment
X5741 N5741 N5742 Segment
X5742 N5742 N5743 Segment
X5743 N5743 N5744 Segment
X5744 N5744 N5745 Segment
X5745 N5745 N5746 Segment
X5746 N5746 N5747 Segment
X5747 N5747 N5748 Segment
X5748 N5748 N5749 Segment
X5749 N5749 N5750 Segment
X5750 N5750 N5751 Segment
X5751 N5751 N5752 Segment
X5752 N5752 N5753 Segment
X5753 N5753 N5754 Segment
X5754 N5754 N5755 Segment
X5755 N5755 N5756 Segment
X5756 N5756 N5757 Segment
X5757 N5757 N5758 Segment
X5758 N5758 N5759 Segment
X5759 N5759 N5760 Segment
X5760 N5760 N5761 Segment
X5761 N5761 N5762 Segment
X5762 N5762 N5763 Segment
X5763 N5763 N5764 Segment
X5764 N5764 N5765 Segment
X5765 N5765 N5766 Segment
X5766 N5766 N5767 Segment
X5767 N5767 N5768 Segment
X5768 N5768 N5769 Segment
X5769 N5769 N5770 Segment
X5770 N5770 N5771 Segment
X5771 N5771 N5772 Segment
X5772 N5772 N5773 Segment
X5773 N5773 N5774 Segment
X5774 N5774 N5775 Segment
X5775 N5775 N5776 Segment
X5776 N5776 N5777 Segment
X5777 N5777 N5778 Segment
X5778 N5778 N5779 Segment
X5779 N5779 N5780 Segment
X5780 N5780 N5781 Segment
X5781 N5781 N5782 Segment
X5782 N5782 N5783 Segment
X5783 N5783 N5784 Segment
X5784 N5784 N5785 Segment
X5785 N5785 N5786 Segment
X5786 N5786 N5787 Segment
X5787 N5787 N5788 Segment
X5788 N5788 N5789 Segment
X5789 N5789 N5790 Segment
X5790 N5790 N5791 Segment
X5791 N5791 N5792 Segment
X5792 N5792 N5793 Segment
X5793 N5793 N5794 Segment
X5794 N5794 N5795 Segment
X5795 N5795 N5796 Segment
X5796 N5796 N5797 Segment
X5797 N5797 N5798 Segment
X5798 N5798 N5799 Segment
X5799 N5799 N5800 Segment
X5800 N5800 N5801 Segment
X5801 N5801 N5802 Segment
X5802 N5802 N5803 Segment
X5803 N5803 N5804 Segment
X5804 N5804 N5805 Segment
X5805 N5805 N5806 Segment
X5806 N5806 N5807 Segment
X5807 N5807 N5808 Segment
X5808 N5808 N5809 Segment
X5809 N5809 N5810 Segment
X5810 N5810 N5811 Segment
X5811 N5811 N5812 Segment
X5812 N5812 N5813 Segment
X5813 N5813 N5814 Segment
X5814 N5814 N5815 Segment
X5815 N5815 N5816 Segment
X5816 N5816 N5817 Segment
X5817 N5817 N5818 Segment
X5818 N5818 N5819 Segment
X5819 N5819 N5820 Segment
X5820 N5820 N5821 Segment
X5821 N5821 N5822 Segment
X5822 N5822 N5823 Segment
X5823 N5823 N5824 Segment
X5824 N5824 N5825 Segment
X5825 N5825 N5826 Segment
X5826 N5826 N5827 Segment
X5827 N5827 N5828 Segment
X5828 N5828 N5829 Segment
X5829 N5829 N5830 Segment
X5830 N5830 N5831 Segment
X5831 N5831 N5832 Segment
X5832 N5832 N5833 Segment
X5833 N5833 N5834 Segment
X5834 N5834 N5835 Segment
X5835 N5835 N5836 Segment
X5836 N5836 N5837 Segment
X5837 N5837 N5838 Segment
X5838 N5838 N5839 Segment
X5839 N5839 N5840 Segment
X5840 N5840 N5841 Segment
X5841 N5841 N5842 Segment
X5842 N5842 N5843 Segment
X5843 N5843 N5844 Segment
X5844 N5844 N5845 Segment
X5845 N5845 N5846 Segment
X5846 N5846 N5847 Segment
X5847 N5847 N5848 Segment
X5848 N5848 N5849 Segment
X5849 N5849 N5850 Segment
X5850 N5850 N5851 Segment
X5851 N5851 N5852 Segment
X5852 N5852 N5853 Segment
X5853 N5853 N5854 Segment
X5854 N5854 N5855 Segment
X5855 N5855 N5856 Segment
X5856 N5856 N5857 Segment
X5857 N5857 N5858 Segment
X5858 N5858 N5859 Segment
X5859 N5859 N5860 Segment
X5860 N5860 N5861 Segment
X5861 N5861 N5862 Segment
X5862 N5862 N5863 Segment
X5863 N5863 N5864 Segment
X5864 N5864 N5865 Segment
X5865 N5865 N5866 Segment
X5866 N5866 N5867 Segment
X5867 N5867 N5868 Segment
X5868 N5868 N5869 Segment
X5869 N5869 N5870 Segment
X5870 N5870 N5871 Segment
X5871 N5871 N5872 Segment
X5872 N5872 N5873 Segment
X5873 N5873 N5874 Segment
X5874 N5874 N5875 Segment
X5875 N5875 N5876 Segment
X5876 N5876 N5877 Segment
X5877 N5877 N5878 Segment
X5878 N5878 N5879 Segment
X5879 N5879 N5880 Segment
X5880 N5880 N5881 Segment
X5881 N5881 N5882 Segment
X5882 N5882 N5883 Segment
X5883 N5883 N5884 Segment
X5884 N5884 N5885 Segment
X5885 N5885 N5886 Segment
X5886 N5886 N5887 Segment
X5887 N5887 N5888 Segment
X5888 N5888 N5889 Segment
X5889 N5889 N5890 Segment
X5890 N5890 N5891 Segment
X5891 N5891 N5892 Segment
X5892 N5892 N5893 Segment
X5893 N5893 N5894 Segment
X5894 N5894 N5895 Segment
X5895 N5895 N5896 Segment
X5896 N5896 N5897 Segment
X5897 N5897 N5898 Segment
X5898 N5898 N5899 Segment
X5899 N5899 N5900 Segment
X5900 N5900 N5901 Segment
X5901 N5901 N5902 Segment
X5902 N5902 N5903 Segment
X5903 N5903 N5904 Segment
X5904 N5904 N5905 Segment
X5905 N5905 N5906 Segment
X5906 N5906 N5907 Segment
X5907 N5907 N5908 Segment
X5908 N5908 N5909 Segment
X5909 N5909 N5910 Segment
X5910 N5910 N5911 Segment
X5911 N5911 N5912 Segment
X5912 N5912 N5913 Segment
X5913 N5913 N5914 Segment
X5914 N5914 N5915 Segment
X5915 N5915 N5916 Segment
X5916 N5916 N5917 Segment
X5917 N5917 N5918 Segment
X5918 N5918 N5919 Segment
X5919 N5919 N5920 Segment
X5920 N5920 N5921 Segment
X5921 N5921 N5922 Segment
X5922 N5922 N5923 Segment
X5923 N5923 N5924 Segment
X5924 N5924 N5925 Segment
X5925 N5925 N5926 Segment
X5926 N5926 N5927 Segment
X5927 N5927 N5928 Segment
X5928 N5928 N5929 Segment
X5929 N5929 N5930 Segment
X5930 N5930 N5931 Segment
X5931 N5931 N5932 Segment
X5932 N5932 N5933 Segment
X5933 N5933 N5934 Segment
X5934 N5934 N5935 Segment
X5935 N5935 N5936 Segment
X5936 N5936 N5937 Segment
X5937 N5937 N5938 Segment
X5938 N5938 N5939 Segment
X5939 N5939 N5940 Segment
X5940 N5940 N5941 Segment
X5941 N5941 N5942 Segment
X5942 N5942 N5943 Segment
X5943 N5943 N5944 Segment
X5944 N5944 N5945 Segment
X5945 N5945 N5946 Segment
X5946 N5946 N5947 Segment
X5947 N5947 N5948 Segment
X5948 N5948 N5949 Segment
X5949 N5949 N5950 Segment
X5950 N5950 N5951 Segment
X5951 N5951 N5952 Segment
X5952 N5952 N5953 Segment
X5953 N5953 N5954 Segment
X5954 N5954 N5955 Segment
X5955 N5955 N5956 Segment
X5956 N5956 N5957 Segment
X5957 N5957 N5958 Segment
X5958 N5958 N5959 Segment
X5959 N5959 N5960 Segment
X5960 N5960 N5961 Segment
X5961 N5961 N5962 Segment
X5962 N5962 N5963 Segment
X5963 N5963 N5964 Segment
X5964 N5964 N5965 Segment
X5965 N5965 N5966 Segment
X5966 N5966 N5967 Segment
X5967 N5967 N5968 Segment
X5968 N5968 N5969 Segment
X5969 N5969 N5970 Segment
X5970 N5970 N5971 Segment
X5971 N5971 N5972 Segment
X5972 N5972 N5973 Segment
X5973 N5973 N5974 Segment
X5974 N5974 N5975 Segment
X5975 N5975 N5976 Segment
X5976 N5976 N5977 Segment
X5977 N5977 N5978 Segment
X5978 N5978 N5979 Segment
X5979 N5979 N5980 Segment
X5980 N5980 N5981 Segment
X5981 N5981 N5982 Segment
X5982 N5982 N5983 Segment
X5983 N5983 N5984 Segment
X5984 N5984 N5985 Segment
X5985 N5985 N5986 Segment
X5986 N5986 N5987 Segment
X5987 N5987 N5988 Segment
X5988 N5988 N5989 Segment
X5989 N5989 N5990 Segment
X5990 N5990 N5991 Segment
X5991 N5991 N5992 Segment
X5992 N5992 N5993 Segment
X5993 N5993 N5994 Segment
X5994 N5994 N5995 Segment
X5995 N5995 N5996 Segment
X5996 N5996 N5997 Segment
X5997 N5997 N5998 Segment
X5998 N5998 N5999 Segment
X5999 N5999 N6000 Segment
X6000 N6000 N6001 Segment
X6001 N6001 N6002 Segment
X6002 N6002 N6003 Segment
X6003 N6003 N6004 Segment
X6004 N6004 N6005 Segment
X6005 N6005 N6006 Segment
X6006 N6006 N6007 Segment
X6007 N6007 N6008 Segment
X6008 N6008 N6009 Segment
X6009 N6009 N6010 Segment
X6010 N6010 N6011 Segment
X6011 N6011 N6012 Segment
X6012 N6012 N6013 Segment
X6013 N6013 N6014 Segment
X6014 N6014 N6015 Segment
X6015 N6015 N6016 Segment
X6016 N6016 N6017 Segment
X6017 N6017 N6018 Segment
X6018 N6018 N6019 Segment
X6019 N6019 N6020 Segment
X6020 N6020 N6021 Segment
X6021 N6021 N6022 Segment
X6022 N6022 N6023 Segment
X6023 N6023 N6024 Segment
X6024 N6024 N6025 Segment
X6025 N6025 N6026 Segment
X6026 N6026 N6027 Segment
X6027 N6027 N6028 Segment
X6028 N6028 N6029 Segment
X6029 N6029 N6030 Segment
X6030 N6030 N6031 Segment
X6031 N6031 N6032 Segment
X6032 N6032 N6033 Segment
X6033 N6033 N6034 Segment
X6034 N6034 N6035 Segment
X6035 N6035 N6036 Segment
X6036 N6036 N6037 Segment
X6037 N6037 N6038 Segment
X6038 N6038 N6039 Segment
X6039 N6039 N6040 Segment
X6040 N6040 N6041 Segment
X6041 N6041 N6042 Segment
X6042 N6042 N6043 Segment
X6043 N6043 N6044 Segment
X6044 N6044 N6045 Segment
X6045 N6045 N6046 Segment
X6046 N6046 N6047 Segment
X6047 N6047 N6048 Segment
X6048 N6048 N6049 Segment
X6049 N6049 N6050 Segment
X6050 N6050 N6051 Segment
X6051 N6051 N6052 Segment
X6052 N6052 N6053 Segment
X6053 N6053 N6054 Segment
X6054 N6054 N6055 Segment
X6055 N6055 N6056 Segment
X6056 N6056 N6057 Segment
X6057 N6057 N6058 Segment
X6058 N6058 N6059 Segment
X6059 N6059 N6060 Segment
X6060 N6060 N6061 Segment
X6061 N6061 N6062 Segment
X6062 N6062 N6063 Segment
X6063 N6063 N6064 Segment
X6064 N6064 N6065 Segment
X6065 N6065 N6066 Segment
X6066 N6066 N6067 Segment
X6067 N6067 N6068 Segment
X6068 N6068 N6069 Segment
X6069 N6069 N6070 Segment
X6070 N6070 N6071 Segment
X6071 N6071 N6072 Segment
X6072 N6072 N6073 Segment
X6073 N6073 N6074 Segment
X6074 N6074 N6075 Segment
X6075 N6075 N6076 Segment
X6076 N6076 N6077 Segment
X6077 N6077 N6078 Segment
X6078 N6078 N6079 Segment
X6079 N6079 N6080 Segment
X6080 N6080 N6081 Segment
X6081 N6081 N6082 Segment
X6082 N6082 N6083 Segment
X6083 N6083 N6084 Segment
X6084 N6084 N6085 Segment
X6085 N6085 N6086 Segment
X6086 N6086 N6087 Segment
X6087 N6087 N6088 Segment
X6088 N6088 N6089 Segment
X6089 N6089 N6090 Segment
X6090 N6090 N6091 Segment
X6091 N6091 N6092 Segment
X6092 N6092 N6093 Segment
X6093 N6093 N6094 Segment
X6094 N6094 N6095 Segment
X6095 N6095 N6096 Segment
X6096 N6096 N6097 Segment
X6097 N6097 N6098 Segment
X6098 N6098 N6099 Segment
X6099 N6099 N6100 Segment
X6100 N6100 N6101 Segment
X6101 N6101 N6102 Segment
X6102 N6102 N6103 Segment
X6103 N6103 N6104 Segment
X6104 N6104 N6105 Segment
X6105 N6105 N6106 Segment
X6106 N6106 N6107 Segment
X6107 N6107 N6108 Segment
X6108 N6108 N6109 Segment
X6109 N6109 N6110 Segment
X6110 N6110 N6111 Segment
X6111 N6111 N6112 Segment
X6112 N6112 N6113 Segment
X6113 N6113 N6114 Segment
X6114 N6114 N6115 Segment
X6115 N6115 N6116 Segment
X6116 N6116 N6117 Segment
X6117 N6117 N6118 Segment
X6118 N6118 N6119 Segment
X6119 N6119 N6120 Segment
X6120 N6120 N6121 Segment
X6121 N6121 N6122 Segment
X6122 N6122 N6123 Segment
X6123 N6123 N6124 Segment
X6124 N6124 N6125 Segment
X6125 N6125 N6126 Segment
X6126 N6126 N6127 Segment
X6127 N6127 N6128 Segment
X6128 N6128 N6129 Segment
X6129 N6129 N6130 Segment
X6130 N6130 N6131 Segment
X6131 N6131 N6132 Segment
X6132 N6132 N6133 Segment
X6133 N6133 N6134 Segment
X6134 N6134 N6135 Segment
X6135 N6135 N6136 Segment
X6136 N6136 N6137 Segment
X6137 N6137 N6138 Segment
X6138 N6138 N6139 Segment
X6139 N6139 N6140 Segment
X6140 N6140 N6141 Segment
X6141 N6141 N6142 Segment
X6142 N6142 N6143 Segment
X6143 N6143 N6144 Segment
X6144 N6144 N6145 Segment
X6145 N6145 N6146 Segment
X6146 N6146 N6147 Segment
X6147 N6147 N6148 Segment
X6148 N6148 N6149 Segment
X6149 N6149 N6150 Segment
X6150 N6150 N6151 Segment
X6151 N6151 N6152 Segment
X6152 N6152 N6153 Segment
X6153 N6153 N6154 Segment
X6154 N6154 N6155 Segment
X6155 N6155 N6156 Segment
X6156 N6156 N6157 Segment
X6157 N6157 N6158 Segment
X6158 N6158 N6159 Segment
X6159 N6159 N6160 Segment
X6160 N6160 N6161 Segment
X6161 N6161 N6162 Segment
X6162 N6162 N6163 Segment
X6163 N6163 N6164 Segment
X6164 N6164 N6165 Segment
X6165 N6165 N6166 Segment
X6166 N6166 N6167 Segment
X6167 N6167 N6168 Segment
X6168 N6168 N6169 Segment
X6169 N6169 N6170 Segment
X6170 N6170 N6171 Segment
X6171 N6171 N6172 Segment
X6172 N6172 N6173 Segment
X6173 N6173 N6174 Segment
X6174 N6174 N6175 Segment
X6175 N6175 N6176 Segment
X6176 N6176 N6177 Segment
X6177 N6177 N6178 Segment
X6178 N6178 N6179 Segment
X6179 N6179 N6180 Segment
X6180 N6180 N6181 Segment
X6181 N6181 N6182 Segment
X6182 N6182 N6183 Segment
X6183 N6183 N6184 Segment
X6184 N6184 N6185 Segment
X6185 N6185 N6186 Segment
X6186 N6186 N6187 Segment
X6187 N6187 N6188 Segment
X6188 N6188 N6189 Segment
X6189 N6189 N6190 Segment
X6190 N6190 N6191 Segment
X6191 N6191 N6192 Segment
X6192 N6192 N6193 Segment
X6193 N6193 N6194 Segment
X6194 N6194 N6195 Segment
X6195 N6195 N6196 Segment
X6196 N6196 N6197 Segment
X6197 N6197 N6198 Segment
X6198 N6198 N6199 Segment
X6199 N6199 N6200 Segment
X6200 N6200 N6201 Segment
X6201 N6201 N6202 Segment
X6202 N6202 N6203 Segment
X6203 N6203 N6204 Segment
X6204 N6204 N6205 Segment
X6205 N6205 N6206 Segment
X6206 N6206 N6207 Segment
X6207 N6207 N6208 Segment
X6208 N6208 N6209 Segment
X6209 N6209 N6210 Segment
X6210 N6210 N6211 Segment
X6211 N6211 N6212 Segment
X6212 N6212 N6213 Segment
X6213 N6213 N6214 Segment
X6214 N6214 N6215 Segment
X6215 N6215 N6216 Segment
X6216 N6216 N6217 Segment
X6217 N6217 N6218 Segment
X6218 N6218 N6219 Segment
X6219 N6219 N6220 Segment
X6220 N6220 N6221 Segment
X6221 N6221 N6222 Segment
X6222 N6222 N6223 Segment
X6223 N6223 N6224 Segment
X6224 N6224 N6225 Segment
X6225 N6225 N6226 Segment
X6226 N6226 N6227 Segment
X6227 N6227 N6228 Segment
X6228 N6228 N6229 Segment
X6229 N6229 N6230 Segment
X6230 N6230 N6231 Segment
X6231 N6231 N6232 Segment
X6232 N6232 N6233 Segment
X6233 N6233 N6234 Segment
X6234 N6234 N6235 Segment
X6235 N6235 N6236 Segment
X6236 N6236 N6237 Segment
X6237 N6237 N6238 Segment
X6238 N6238 N6239 Segment
X6239 N6239 N6240 Segment
X6240 N6240 N6241 Segment
X6241 N6241 N6242 Segment
X6242 N6242 N6243 Segment
X6243 N6243 N6244 Segment
X6244 N6244 N6245 Segment
X6245 N6245 N6246 Segment
X6246 N6246 N6247 Segment
X6247 N6247 N6248 Segment
X6248 N6248 N6249 Segment
X6249 N6249 N6250 Segment
X6250 N6250 N6251 Segment
X6251 N6251 N6252 Segment
X6252 N6252 N6253 Segment
X6253 N6253 N6254 Segment
X6254 N6254 N6255 Segment
X6255 N6255 N6256 Segment
X6256 N6256 N6257 Segment
X6257 N6257 N6258 Segment
X6258 N6258 N6259 Segment
X6259 N6259 N6260 Segment
X6260 N6260 N6261 Segment
X6261 N6261 N6262 Segment
X6262 N6262 N6263 Segment
X6263 N6263 N6264 Segment
X6264 N6264 N6265 Segment
X6265 N6265 N6266 Segment
X6266 N6266 N6267 Segment
X6267 N6267 N6268 Segment
X6268 N6268 N6269 Segment
X6269 N6269 N6270 Segment
X6270 N6270 N6271 Segment
X6271 N6271 N6272 Segment
X6272 N6272 N6273 Segment
X6273 N6273 N6274 Segment
X6274 N6274 N6275 Segment
X6275 N6275 N6276 Segment
X6276 N6276 N6277 Segment
X6277 N6277 N6278 Segment
X6278 N6278 N6279 Segment
X6279 N6279 N6280 Segment
X6280 N6280 N6281 Segment
X6281 N6281 N6282 Segment
X6282 N6282 N6283 Segment
X6283 N6283 N6284 Segment
X6284 N6284 N6285 Segment
X6285 N6285 N6286 Segment
X6286 N6286 N6287 Segment
X6287 N6287 N6288 Segment
X6288 N6288 N6289 Segment
X6289 N6289 N6290 Segment
X6290 N6290 N6291 Segment
X6291 N6291 N6292 Segment
X6292 N6292 N6293 Segment
X6293 N6293 N6294 Segment
X6294 N6294 N6295 Segment
X6295 N6295 N6296 Segment
X6296 N6296 N6297 Segment
X6297 N6297 N6298 Segment
X6298 N6298 N6299 Segment
X6299 N6299 N6300 Segment
X6300 N6300 N6301 Segment
X6301 N6301 N6302 Segment
X6302 N6302 N6303 Segment
X6303 N6303 N6304 Segment
X6304 N6304 N6305 Segment
X6305 N6305 N6306 Segment
X6306 N6306 N6307 Segment
X6307 N6307 N6308 Segment
X6308 N6308 N6309 Segment
X6309 N6309 N6310 Segment
X6310 N6310 N6311 Segment
X6311 N6311 N6312 Segment
X6312 N6312 N6313 Segment
X6313 N6313 N6314 Segment
X6314 N6314 N6315 Segment
X6315 N6315 N6316 Segment
X6316 N6316 N6317 Segment
X6317 N6317 N6318 Segment
X6318 N6318 N6319 Segment
X6319 N6319 N6320 Segment
X6320 N6320 N6321 Segment
X6321 N6321 N6322 Segment
X6322 N6322 N6323 Segment
X6323 N6323 N6324 Segment
X6324 N6324 N6325 Segment
X6325 N6325 N6326 Segment
X6326 N6326 N6327 Segment
X6327 N6327 N6328 Segment
X6328 N6328 N6329 Segment
X6329 N6329 N6330 Segment
X6330 N6330 N6331 Segment
X6331 N6331 N6332 Segment
X6332 N6332 N6333 Segment
X6333 N6333 N6334 Segment
X6334 N6334 N6335 Segment
X6335 N6335 N6336 Segment
X6336 N6336 N6337 Segment
X6337 N6337 N6338 Segment
X6338 N6338 N6339 Segment
X6339 N6339 N6340 Segment
X6340 N6340 N6341 Segment
X6341 N6341 N6342 Segment
X6342 N6342 N6343 Segment
X6343 N6343 N6344 Segment
X6344 N6344 N6345 Segment
X6345 N6345 N6346 Segment
X6346 N6346 N6347 Segment
X6347 N6347 N6348 Segment
X6348 N6348 N6349 Segment
X6349 N6349 N6350 Segment
X6350 N6350 N6351 Segment
X6351 N6351 N6352 Segment
X6352 N6352 N6353 Segment
X6353 N6353 N6354 Segment
X6354 N6354 N6355 Segment
X6355 N6355 N6356 Segment
X6356 N6356 N6357 Segment
X6357 N6357 N6358 Segment
X6358 N6358 N6359 Segment
X6359 N6359 N6360 Segment
X6360 N6360 N6361 Segment
X6361 N6361 N6362 Segment
X6362 N6362 N6363 Segment
X6363 N6363 N6364 Segment
X6364 N6364 N6365 Segment
X6365 N6365 N6366 Segment
X6366 N6366 N6367 Segment
X6367 N6367 N6368 Segment
X6368 N6368 N6369 Segment
X6369 N6369 N6370 Segment
X6370 N6370 N6371 Segment
X6371 N6371 N6372 Segment
X6372 N6372 N6373 Segment
X6373 N6373 N6374 Segment
X6374 N6374 N6375 Segment
X6375 N6375 N6376 Segment
X6376 N6376 N6377 Segment
X6377 N6377 N6378 Segment
X6378 N6378 N6379 Segment
X6379 N6379 N6380 Segment
X6380 N6380 N6381 Segment
X6381 N6381 N6382 Segment
X6382 N6382 N6383 Segment
X6383 N6383 N6384 Segment
X6384 N6384 N6385 Segment
X6385 N6385 N6386 Segment
X6386 N6386 N6387 Segment
X6387 N6387 N6388 Segment
X6388 N6388 N6389 Segment
X6389 N6389 N6390 Segment
X6390 N6390 N6391 Segment
X6391 N6391 N6392 Segment
X6392 N6392 N6393 Segment
X6393 N6393 N6394 Segment
X6394 N6394 N6395 Segment
X6395 N6395 N6396 Segment
X6396 N6396 N6397 Segment
X6397 N6397 N6398 Segment
X6398 N6398 N6399 Segment
X6399 N6399 N6400 Segment
X6400 N6400 N6401 Segment
X6401 N6401 N6402 Segment
X6402 N6402 N6403 Segment
X6403 N6403 N6404 Segment
X6404 N6404 N6405 Segment
X6405 N6405 N6406 Segment
X6406 N6406 N6407 Segment
X6407 N6407 N6408 Segment
X6408 N6408 N6409 Segment
X6409 N6409 N6410 Segment
X6410 N6410 N6411 Segment
X6411 N6411 N6412 Segment
X6412 N6412 N6413 Segment
X6413 N6413 N6414 Segment
X6414 N6414 N6415 Segment
X6415 N6415 N6416 Segment
X6416 N6416 N6417 Segment
X6417 N6417 N6418 Segment
X6418 N6418 N6419 Segment
X6419 N6419 N6420 Segment
X6420 N6420 N6421 Segment
X6421 N6421 N6422 Segment
X6422 N6422 N6423 Segment
X6423 N6423 N6424 Segment
X6424 N6424 N6425 Segment
X6425 N6425 N6426 Segment
X6426 N6426 N6427 Segment
X6427 N6427 N6428 Segment
X6428 N6428 N6429 Segment
X6429 N6429 N6430 Segment
X6430 N6430 N6431 Segment
X6431 N6431 N6432 Segment
X6432 N6432 N6433 Segment
X6433 N6433 N6434 Segment
X6434 N6434 N6435 Segment
X6435 N6435 N6436 Segment
X6436 N6436 N6437 Segment
X6437 N6437 N6438 Segment
X6438 N6438 N6439 Segment
X6439 N6439 N6440 Segment
X6440 N6440 N6441 Segment
X6441 N6441 N6442 Segment
X6442 N6442 N6443 Segment
X6443 N6443 N6444 Segment
X6444 N6444 N6445 Segment
X6445 N6445 N6446 Segment
X6446 N6446 N6447 Segment
X6447 N6447 N6448 Segment
X6448 N6448 N6449 Segment
X6449 N6449 N6450 Segment
X6450 N6450 N6451 Segment
X6451 N6451 N6452 Segment
X6452 N6452 N6453 Segment
X6453 N6453 N6454 Segment
X6454 N6454 N6455 Segment
X6455 N6455 N6456 Segment
X6456 N6456 N6457 Segment
X6457 N6457 N6458 Segment
X6458 N6458 N6459 Segment
X6459 N6459 N6460 Segment
X6460 N6460 N6461 Segment
X6461 N6461 N6462 Segment
X6462 N6462 N6463 Segment
X6463 N6463 N6464 Segment
X6464 N6464 N6465 Segment
X6465 N6465 N6466 Segment
X6466 N6466 N6467 Segment
X6467 N6467 N6468 Segment
X6468 N6468 N6469 Segment
X6469 N6469 N6470 Segment
X6470 N6470 N6471 Segment
X6471 N6471 N6472 Segment
X6472 N6472 N6473 Segment
X6473 N6473 N6474 Segment
X6474 N6474 N6475 Segment
X6475 N6475 N6476 Segment
X6476 N6476 N6477 Segment
X6477 N6477 N6478 Segment
X6478 N6478 N6479 Segment
X6479 N6479 N6480 Segment
X6480 N6480 N6481 Segment
X6481 N6481 N6482 Segment
X6482 N6482 N6483 Segment
X6483 N6483 N6484 Segment
X6484 N6484 N6485 Segment
X6485 N6485 N6486 Segment
X6486 N6486 N6487 Segment
X6487 N6487 N6488 Segment
X6488 N6488 N6489 Segment
X6489 N6489 N6490 Segment
X6490 N6490 N6491 Segment
X6491 N6491 N6492 Segment
X6492 N6492 N6493 Segment
X6493 N6493 N6494 Segment
X6494 N6494 N6495 Segment
X6495 N6495 N6496 Segment
X6496 N6496 N6497 Segment
X6497 N6497 N6498 Segment
X6498 N6498 N6499 Segment
X6499 N6499 N6500 Segment
X6500 N6500 N6501 Segment
X6501 N6501 N6502 Segment
X6502 N6502 N6503 Segment
X6503 N6503 N6504 Segment
X6504 N6504 N6505 Segment
X6505 N6505 N6506 Segment
X6506 N6506 N6507 Segment
X6507 N6507 N6508 Segment
X6508 N6508 N6509 Segment
X6509 N6509 N6510 Segment
X6510 N6510 N6511 Segment
X6511 N6511 N6512 Segment
X6512 N6512 N6513 Segment
X6513 N6513 N6514 Segment
X6514 N6514 N6515 Segment
X6515 N6515 N6516 Segment
X6516 N6516 N6517 Segment
X6517 N6517 N6518 Segment
X6518 N6518 N6519 Segment
X6519 N6519 N6520 Segment
X6520 N6520 N6521 Segment
X6521 N6521 N6522 Segment
X6522 N6522 N6523 Segment
X6523 N6523 N6524 Segment
X6524 N6524 N6525 Segment
X6525 N6525 N6526 Segment
X6526 N6526 N6527 Segment
X6527 N6527 N6528 Segment
X6528 N6528 N6529 Segment
X6529 N6529 N6530 Segment
X6530 N6530 N6531 Segment
X6531 N6531 N6532 Segment
X6532 N6532 N6533 Segment
X6533 N6533 N6534 Segment
X6534 N6534 N6535 Segment
X6535 N6535 N6536 Segment
X6536 N6536 N6537 Segment
X6537 N6537 N6538 Segment
X6538 N6538 N6539 Segment
X6539 N6539 N6540 Segment
X6540 N6540 N6541 Segment
X6541 N6541 N6542 Segment
X6542 N6542 N6543 Segment
X6543 N6543 N6544 Segment
X6544 N6544 N6545 Segment
X6545 N6545 N6546 Segment
X6546 N6546 N6547 Segment
X6547 N6547 N6548 Segment
X6548 N6548 N6549 Segment
X6549 N6549 N6550 Segment
X6550 N6550 N6551 Segment
X6551 N6551 N6552 Segment
X6552 N6552 N6553 Segment
X6553 N6553 N6554 Segment
X6554 N6554 N6555 Segment
X6555 N6555 N6556 Segment
X6556 N6556 N6557 Segment
X6557 N6557 N6558 Segment
X6558 N6558 N6559 Segment
X6559 N6559 N6560 Segment
X6560 N6560 N6561 Segment
X6561 N6561 N6562 Segment
X6562 N6562 N6563 Segment
X6563 N6563 N6564 Segment
X6564 N6564 N6565 Segment
X6565 N6565 N6566 Segment
X6566 N6566 N6567 Segment
X6567 N6567 N6568 Segment
X6568 N6568 N6569 Segment
X6569 N6569 N6570 Segment
X6570 N6570 N6571 Segment
X6571 N6571 N6572 Segment
X6572 N6572 N6573 Segment
X6573 N6573 N6574 Segment
X6574 N6574 N6575 Segment
X6575 N6575 N6576 Segment
X6576 N6576 N6577 Segment
X6577 N6577 N6578 Segment
X6578 N6578 N6579 Segment
X6579 N6579 N6580 Segment
X6580 N6580 N6581 Segment
X6581 N6581 N6582 Segment
X6582 N6582 N6583 Segment
X6583 N6583 N6584 Segment
X6584 N6584 N6585 Segment
X6585 N6585 N6586 Segment
X6586 N6586 N6587 Segment
X6587 N6587 N6588 Segment
X6588 N6588 N6589 Segment
X6589 N6589 N6590 Segment
X6590 N6590 N6591 Segment
X6591 N6591 N6592 Segment
X6592 N6592 N6593 Segment
X6593 N6593 N6594 Segment
X6594 N6594 N6595 Segment
X6595 N6595 N6596 Segment
X6596 N6596 N6597 Segment
X6597 N6597 N6598 Segment
X6598 N6598 N6599 Segment
X6599 N6599 N6600 Segment
X6600 N6600 N6601 Segment
X6601 N6601 N6602 Segment
X6602 N6602 N6603 Segment
X6603 N6603 N6604 Segment
X6604 N6604 N6605 Segment
X6605 N6605 N6606 Segment
X6606 N6606 N6607 Segment
X6607 N6607 N6608 Segment
X6608 N6608 N6609 Segment
X6609 N6609 N6610 Segment
X6610 N6610 N6611 Segment
X6611 N6611 N6612 Segment
X6612 N6612 N6613 Segment
X6613 N6613 N6614 Segment
X6614 N6614 N6615 Segment
X6615 N6615 N6616 Segment
X6616 N6616 N6617 Segment
X6617 N6617 N6618 Segment
X6618 N6618 N6619 Segment
X6619 N6619 N6620 Segment
X6620 N6620 N6621 Segment
X6621 N6621 N6622 Segment
X6622 N6622 N6623 Segment
X6623 N6623 N6624 Segment
X6624 N6624 N6625 Segment
X6625 N6625 N6626 Segment
X6626 N6626 N6627 Segment
X6627 N6627 N6628 Segment
X6628 N6628 N6629 Segment
X6629 N6629 N6630 Segment
X6630 N6630 N6631 Segment
X6631 N6631 N6632 Segment
X6632 N6632 N6633 Segment
X6633 N6633 N6634 Segment
X6634 N6634 N6635 Segment
X6635 N6635 N6636 Segment
X6636 N6636 N6637 Segment
X6637 N6637 N6638 Segment
X6638 N6638 N6639 Segment
X6639 N6639 N6640 Segment
X6640 N6640 N6641 Segment
X6641 N6641 N6642 Segment
X6642 N6642 N6643 Segment
X6643 N6643 N6644 Segment
X6644 N6644 N6645 Segment
X6645 N6645 N6646 Segment
X6646 N6646 N6647 Segment
X6647 N6647 N6648 Segment
X6648 N6648 N6649 Segment
X6649 N6649 N6650 Segment
X6650 N6650 N6651 Segment
X6651 N6651 N6652 Segment
X6652 N6652 N6653 Segment
X6653 N6653 N6654 Segment
X6654 N6654 N6655 Segment
X6655 N6655 N6656 Segment
X6656 N6656 N6657 Segment
X6657 N6657 N6658 Segment
X6658 N6658 N6659 Segment
X6659 N6659 N6660 Segment
X6660 N6660 N6661 Segment
X6661 N6661 N6662 Segment
X6662 N6662 N6663 Segment
X6663 N6663 N6664 Segment
X6664 N6664 N6665 Segment
X6665 N6665 N6666 Segment
X6666 N6666 N6667 Segment
X6667 N6667 N6668 Segment
X6668 N6668 N6669 Segment
X6669 N6669 N6670 Segment
X6670 N6670 N6671 Segment
X6671 N6671 N6672 Segment
X6672 N6672 N6673 Segment
X6673 N6673 N6674 Segment
X6674 N6674 N6675 Segment
X6675 N6675 N6676 Segment
X6676 N6676 N6677 Segment
X6677 N6677 N6678 Segment
X6678 N6678 N6679 Segment
X6679 N6679 N6680 Segment
X6680 N6680 N6681 Segment
X6681 N6681 N6682 Segment
X6682 N6682 N6683 Segment
X6683 N6683 N6684 Segment
X6684 N6684 N6685 Segment
X6685 N6685 N6686 Segment
X6686 N6686 N6687 Segment
X6687 N6687 N6688 Segment
X6688 N6688 N6689 Segment
X6689 N6689 N6690 Segment
X6690 N6690 N6691 Segment
X6691 N6691 N6692 Segment
X6692 N6692 N6693 Segment
X6693 N6693 N6694 Segment
X6694 N6694 N6695 Segment
X6695 N6695 N6696 Segment
X6696 N6696 N6697 Segment
X6697 N6697 N6698 Segment
X6698 N6698 N6699 Segment
X6699 N6699 N6700 Segment
X6700 N6700 N6701 Segment
X6701 N6701 N6702 Segment
X6702 N6702 N6703 Segment
X6703 N6703 N6704 Segment
X6704 N6704 N6705 Segment
X6705 N6705 N6706 Segment
X6706 N6706 N6707 Segment
X6707 N6707 N6708 Segment
X6708 N6708 N6709 Segment
X6709 N6709 N6710 Segment
X6710 N6710 N6711 Segment
X6711 N6711 N6712 Segment
X6712 N6712 N6713 Segment
X6713 N6713 N6714 Segment
X6714 N6714 N6715 Segment
X6715 N6715 N6716 Segment
X6716 N6716 N6717 Segment
X6717 N6717 N6718 Segment
X6718 N6718 N6719 Segment
X6719 N6719 N6720 Segment
X6720 N6720 N6721 Segment
X6721 N6721 N6722 Segment
X6722 N6722 N6723 Segment
X6723 N6723 N6724 Segment
X6724 N6724 N6725 Segment
X6725 N6725 N6726 Segment
X6726 N6726 N6727 Segment
X6727 N6727 N6728 Segment
X6728 N6728 N6729 Segment
X6729 N6729 N6730 Segment
X6730 N6730 N6731 Segment
X6731 N6731 N6732 Segment
X6732 N6732 N6733 Segment
X6733 N6733 N6734 Segment
X6734 N6734 N6735 Segment
X6735 N6735 N6736 Segment
X6736 N6736 N6737 Segment
X6737 N6737 N6738 Segment
X6738 N6738 N6739 Segment
X6739 N6739 N6740 Segment
X6740 N6740 N6741 Segment
X6741 N6741 N6742 Segment
X6742 N6742 N6743 Segment
X6743 N6743 N6744 Segment
X6744 N6744 N6745 Segment
X6745 N6745 N6746 Segment
X6746 N6746 N6747 Segment
X6747 N6747 N6748 Segment
X6748 N6748 N6749 Segment
X6749 N6749 N6750 Segment
X6750 N6750 N6751 Segment
X6751 N6751 N6752 Segment
X6752 N6752 N6753 Segment
X6753 N6753 N6754 Segment
X6754 N6754 N6755 Segment
X6755 N6755 N6756 Segment
X6756 N6756 N6757 Segment
X6757 N6757 N6758 Segment
X6758 N6758 N6759 Segment
X6759 N6759 N6760 Segment
X6760 N6760 N6761 Segment
X6761 N6761 N6762 Segment
X6762 N6762 N6763 Segment
X6763 N6763 N6764 Segment
X6764 N6764 N6765 Segment
X6765 N6765 N6766 Segment
X6766 N6766 N6767 Segment
X6767 N6767 N6768 Segment
X6768 N6768 N6769 Segment
X6769 N6769 N6770 Segment
X6770 N6770 N6771 Segment
X6771 N6771 N6772 Segment
X6772 N6772 N6773 Segment
X6773 N6773 N6774 Segment
X6774 N6774 N6775 Segment
X6775 N6775 N6776 Segment
X6776 N6776 N6777 Segment
X6777 N6777 N6778 Segment
X6778 N6778 N6779 Segment
X6779 N6779 N6780 Segment
X6780 N6780 N6781 Segment
X6781 N6781 N6782 Segment
X6782 N6782 N6783 Segment
X6783 N6783 N6784 Segment
X6784 N6784 N6785 Segment
X6785 N6785 N6786 Segment
X6786 N6786 N6787 Segment
X6787 N6787 N6788 Segment
X6788 N6788 N6789 Segment
X6789 N6789 N6790 Segment
X6790 N6790 N6791 Segment
X6791 N6791 N6792 Segment
X6792 N6792 N6793 Segment
X6793 N6793 N6794 Segment
X6794 N6794 N6795 Segment
X6795 N6795 N6796 Segment
X6796 N6796 N6797 Segment
X6797 N6797 N6798 Segment
X6798 N6798 N6799 Segment
X6799 N6799 N6800 Segment
X6800 N6800 N6801 Segment
X6801 N6801 N6802 Segment
X6802 N6802 N6803 Segment
X6803 N6803 N6804 Segment
X6804 N6804 N6805 Segment
X6805 N6805 N6806 Segment
X6806 N6806 N6807 Segment
X6807 N6807 N6808 Segment
X6808 N6808 N6809 Segment
X6809 N6809 N6810 Segment
X6810 N6810 N6811 Segment
X6811 N6811 N6812 Segment
X6812 N6812 N6813 Segment
X6813 N6813 N6814 Segment
X6814 N6814 N6815 Segment
X6815 N6815 N6816 Segment
X6816 N6816 N6817 Segment
X6817 N6817 N6818 Segment
X6818 N6818 N6819 Segment
X6819 N6819 N6820 Segment
X6820 N6820 N6821 Segment
X6821 N6821 N6822 Segment
X6822 N6822 N6823 Segment
X6823 N6823 N6824 Segment
X6824 N6824 N6825 Segment
X6825 N6825 N6826 Segment
X6826 N6826 N6827 Segment
X6827 N6827 N6828 Segment
X6828 N6828 N6829 Segment
X6829 N6829 N6830 Segment
X6830 N6830 N6831 Segment
X6831 N6831 N6832 Segment
X6832 N6832 N6833 Segment
X6833 N6833 N6834 Segment
X6834 N6834 N6835 Segment
X6835 N6835 N6836 Segment
X6836 N6836 N6837 Segment
X6837 N6837 N6838 Segment
X6838 N6838 N6839 Segment
X6839 N6839 N6840 Segment
X6840 N6840 N6841 Segment
X6841 N6841 N6842 Segment
X6842 N6842 N6843 Segment
X6843 N6843 N6844 Segment
X6844 N6844 N6845 Segment
X6845 N6845 N6846 Segment
X6846 N6846 N6847 Segment
X6847 N6847 N6848 Segment
X6848 N6848 N6849 Segment
X6849 N6849 N6850 Segment
X6850 N6850 N6851 Segment
X6851 N6851 N6852 Segment
X6852 N6852 N6853 Segment
X6853 N6853 N6854 Segment
X6854 N6854 N6855 Segment
X6855 N6855 N6856 Segment
X6856 N6856 N6857 Segment
X6857 N6857 N6858 Segment
X6858 N6858 N6859 Segment
X6859 N6859 N6860 Segment
X6860 N6860 N6861 Segment
X6861 N6861 N6862 Segment
X6862 N6862 N6863 Segment
X6863 N6863 N6864 Segment
X6864 N6864 N6865 Segment
X6865 N6865 N6866 Segment
X6866 N6866 N6867 Segment
X6867 N6867 N6868 Segment
X6868 N6868 N6869 Segment
X6869 N6869 N6870 Segment
X6870 N6870 N6871 Segment
X6871 N6871 N6872 Segment
X6872 N6872 N6873 Segment
X6873 N6873 N6874 Segment
X6874 N6874 N6875 Segment
X6875 N6875 N6876 Segment
X6876 N6876 N6877 Segment
X6877 N6877 N6878 Segment
X6878 N6878 N6879 Segment
X6879 N6879 N6880 Segment
X6880 N6880 N6881 Segment
X6881 N6881 N6882 Segment
X6882 N6882 N6883 Segment
X6883 N6883 N6884 Segment
X6884 N6884 N6885 Segment
X6885 N6885 N6886 Segment
X6886 N6886 N6887 Segment
X6887 N6887 N6888 Segment
X6888 N6888 N6889 Segment
X6889 N6889 N6890 Segment
X6890 N6890 N6891 Segment
X6891 N6891 N6892 Segment
X6892 N6892 N6893 Segment
X6893 N6893 N6894 Segment
X6894 N6894 N6895 Segment
X6895 N6895 N6896 Segment
X6896 N6896 N6897 Segment
X6897 N6897 N6898 Segment
X6898 N6898 N6899 Segment
X6899 N6899 N6900 Segment
X6900 N6900 N6901 Segment
X6901 N6901 N6902 Segment
X6902 N6902 N6903 Segment
X6903 N6903 N6904 Segment
X6904 N6904 N6905 Segment
X6905 N6905 N6906 Segment
X6906 N6906 N6907 Segment
X6907 N6907 N6908 Segment
X6908 N6908 N6909 Segment
X6909 N6909 N6910 Segment
X6910 N6910 N6911 Segment
X6911 N6911 N6912 Segment
X6912 N6912 N6913 Segment
X6913 N6913 N6914 Segment
X6914 N6914 N6915 Segment
X6915 N6915 N6916 Segment
X6916 N6916 N6917 Segment
X6917 N6917 N6918 Segment
X6918 N6918 N6919 Segment
X6919 N6919 N6920 Segment
X6920 N6920 N6921 Segment
X6921 N6921 N6922 Segment
X6922 N6922 N6923 Segment
X6923 N6923 N6924 Segment
X6924 N6924 N6925 Segment
X6925 N6925 N6926 Segment
X6926 N6926 N6927 Segment
X6927 N6927 N6928 Segment
X6928 N6928 N6929 Segment
X6929 N6929 N6930 Segment
X6930 N6930 N6931 Segment
X6931 N6931 N6932 Segment
X6932 N6932 N6933 Segment
X6933 N6933 N6934 Segment
X6934 N6934 N6935 Segment
X6935 N6935 N6936 Segment
X6936 N6936 N6937 Segment
X6937 N6937 N6938 Segment
X6938 N6938 N6939 Segment
X6939 N6939 N6940 Segment
X6940 N6940 N6941 Segment
X6941 N6941 N6942 Segment
X6942 N6942 N6943 Segment
X6943 N6943 N6944 Segment
X6944 N6944 N6945 Segment
X6945 N6945 N6946 Segment
X6946 N6946 N6947 Segment
X6947 N6947 N6948 Segment
X6948 N6948 N6949 Segment
X6949 N6949 N6950 Segment
X6950 N6950 N6951 Segment
X6951 N6951 N6952 Segment
X6952 N6952 N6953 Segment
X6953 N6953 N6954 Segment
X6954 N6954 N6955 Segment
X6955 N6955 N6956 Segment
X6956 N6956 N6957 Segment
X6957 N6957 N6958 Segment
X6958 N6958 N6959 Segment
X6959 N6959 N6960 Segment
X6960 N6960 N6961 Segment
X6961 N6961 N6962 Segment
X6962 N6962 N6963 Segment
X6963 N6963 N6964 Segment
X6964 N6964 N6965 Segment
X6965 N6965 N6966 Segment
X6966 N6966 N6967 Segment
X6967 N6967 N6968 Segment
X6968 N6968 N6969 Segment
X6969 N6969 N6970 Segment
X6970 N6970 N6971 Segment
X6971 N6971 N6972 Segment
X6972 N6972 N6973 Segment
X6973 N6973 N6974 Segment
X6974 N6974 N6975 Segment
X6975 N6975 N6976 Segment
X6976 N6976 N6977 Segment
X6977 N6977 N6978 Segment
X6978 N6978 N6979 Segment
X6979 N6979 N6980 Segment
X6980 N6980 N6981 Segment
X6981 N6981 N6982 Segment
X6982 N6982 N6983 Segment
X6983 N6983 N6984 Segment
X6984 N6984 N6985 Segment
X6985 N6985 N6986 Segment
X6986 N6986 N6987 Segment
X6987 N6987 N6988 Segment
X6988 N6988 N6989 Segment
X6989 N6989 N6990 Segment
X6990 N6990 N6991 Segment
X6991 N6991 N6992 Segment
X6992 N6992 N6993 Segment
X6993 N6993 N6994 Segment
X6994 N6994 N6995 Segment
X6995 N6995 N6996 Segment
X6996 N6996 N6997 Segment
X6997 N6997 N6998 Segment
X6998 N6998 N6999 Segment
X6999 N6999 N7000 Segment
X7000 N7000 N7001 Segment
X7001 N7001 N7002 Segment
X7002 N7002 N7003 Segment
X7003 N7003 N7004 Segment
X7004 N7004 N7005 Segment
X7005 N7005 N7006 Segment
X7006 N7006 N7007 Segment
X7007 N7007 N7008 Segment
X7008 N7008 N7009 Segment
X7009 N7009 N7010 Segment
X7010 N7010 N7011 Segment
X7011 N7011 N7012 Segment
X7012 N7012 N7013 Segment
X7013 N7013 N7014 Segment
X7014 N7014 N7015 Segment
X7015 N7015 N7016 Segment
X7016 N7016 N7017 Segment
X7017 N7017 N7018 Segment
X7018 N7018 N7019 Segment
X7019 N7019 N7020 Segment
X7020 N7020 N7021 Segment
X7021 N7021 N7022 Segment
X7022 N7022 N7023 Segment
X7023 N7023 N7024 Segment
X7024 N7024 N7025 Segment
X7025 N7025 N7026 Segment
X7026 N7026 N7027 Segment
X7027 N7027 N7028 Segment
X7028 N7028 N7029 Segment
X7029 N7029 N7030 Segment
X7030 N7030 N7031 Segment
X7031 N7031 N7032 Segment
X7032 N7032 N7033 Segment
X7033 N7033 N7034 Segment
X7034 N7034 N7035 Segment
X7035 N7035 N7036 Segment
X7036 N7036 N7037 Segment
X7037 N7037 N7038 Segment
X7038 N7038 N7039 Segment
X7039 N7039 N7040 Segment
X7040 N7040 N7041 Segment
X7041 N7041 N7042 Segment
X7042 N7042 N7043 Segment
X7043 N7043 N7044 Segment
X7044 N7044 N7045 Segment
X7045 N7045 N7046 Segment
X7046 N7046 N7047 Segment
X7047 N7047 N7048 Segment
X7048 N7048 N7049 Segment
X7049 N7049 N7050 Segment
X7050 N7050 N7051 Segment
X7051 N7051 N7052 Segment
X7052 N7052 N7053 Segment
X7053 N7053 N7054 Segment
X7054 N7054 N7055 Segment
X7055 N7055 N7056 Segment
X7056 N7056 N7057 Segment
X7057 N7057 N7058 Segment
X7058 N7058 N7059 Segment
X7059 N7059 N7060 Segment
X7060 N7060 N7061 Segment
X7061 N7061 N7062 Segment
X7062 N7062 N7063 Segment
X7063 N7063 N7064 Segment
X7064 N7064 N7065 Segment
X7065 N7065 N7066 Segment
X7066 N7066 N7067 Segment
X7067 N7067 N7068 Segment
X7068 N7068 N7069 Segment
X7069 N7069 N7070 Segment
X7070 N7070 N7071 Segment
X7071 N7071 N7072 Segment
X7072 N7072 N7073 Segment
X7073 N7073 N7074 Segment
X7074 N7074 N7075 Segment
X7075 N7075 N7076 Segment
X7076 N7076 N7077 Segment
X7077 N7077 N7078 Segment
X7078 N7078 N7079 Segment
X7079 N7079 N7080 Segment
X7080 N7080 N7081 Segment
X7081 N7081 N7082 Segment
X7082 N7082 N7083 Segment
X7083 N7083 N7084 Segment
X7084 N7084 N7085 Segment
X7085 N7085 N7086 Segment
X7086 N7086 N7087 Segment
X7087 N7087 N7088 Segment
X7088 N7088 N7089 Segment
X7089 N7089 N7090 Segment
X7090 N7090 N7091 Segment
X7091 N7091 N7092 Segment
X7092 N7092 N7093 Segment
X7093 N7093 N7094 Segment
X7094 N7094 N7095 Segment
X7095 N7095 N7096 Segment
X7096 N7096 N7097 Segment
X7097 N7097 N7098 Segment
X7098 N7098 N7099 Segment
X7099 N7099 N7100 Segment
X7100 N7100 N7101 Segment
X7101 N7101 N7102 Segment
X7102 N7102 N7103 Segment
X7103 N7103 N7104 Segment
X7104 N7104 N7105 Segment
X7105 N7105 N7106 Segment
X7106 N7106 N7107 Segment
X7107 N7107 N7108 Segment
X7108 N7108 N7109 Segment
X7109 N7109 N7110 Segment
X7110 N7110 N7111 Segment
X7111 N7111 N7112 Segment
X7112 N7112 N7113 Segment
X7113 N7113 N7114 Segment
X7114 N7114 N7115 Segment
X7115 N7115 N7116 Segment
X7116 N7116 N7117 Segment
X7117 N7117 N7118 Segment
X7118 N7118 N7119 Segment
X7119 N7119 N7120 Segment
X7120 N7120 N7121 Segment
X7121 N7121 N7122 Segment
X7122 N7122 N7123 Segment
X7123 N7123 N7124 Segment
X7124 N7124 N7125 Segment
X7125 N7125 N7126 Segment
X7126 N7126 N7127 Segment
X7127 N7127 N7128 Segment
X7128 N7128 N7129 Segment
X7129 N7129 N7130 Segment
X7130 N7130 N7131 Segment
X7131 N7131 N7132 Segment
X7132 N7132 N7133 Segment
X7133 N7133 N7134 Segment
X7134 N7134 N7135 Segment
X7135 N7135 N7136 Segment
X7136 N7136 N7137 Segment
X7137 N7137 N7138 Segment
X7138 N7138 N7139 Segment
X7139 N7139 N7140 Segment
X7140 N7140 N7141 Segment
X7141 N7141 N7142 Segment
X7142 N7142 N7143 Segment
X7143 N7143 N7144 Segment
X7144 N7144 N7145 Segment
X7145 N7145 N7146 Segment
X7146 N7146 N7147 Segment
X7147 N7147 N7148 Segment
X7148 N7148 N7149 Segment
X7149 N7149 N7150 Segment
X7150 N7150 N7151 Segment
X7151 N7151 N7152 Segment
X7152 N7152 N7153 Segment
X7153 N7153 N7154 Segment
X7154 N7154 N7155 Segment
X7155 N7155 N7156 Segment
X7156 N7156 N7157 Segment
X7157 N7157 N7158 Segment
X7158 N7158 N7159 Segment
X7159 N7159 N7160 Segment
X7160 N7160 N7161 Segment
X7161 N7161 N7162 Segment
X7162 N7162 N7163 Segment
X7163 N7163 N7164 Segment
X7164 N7164 N7165 Segment
X7165 N7165 N7166 Segment
X7166 N7166 N7167 Segment
X7167 N7167 N7168 Segment
X7168 N7168 N7169 Segment
X7169 N7169 N7170 Segment
X7170 N7170 N7171 Segment
X7171 N7171 N7172 Segment
X7172 N7172 N7173 Segment
X7173 N7173 N7174 Segment
X7174 N7174 N7175 Segment
X7175 N7175 N7176 Segment
X7176 N7176 N7177 Segment
X7177 N7177 N7178 Segment
X7178 N7178 N7179 Segment
X7179 N7179 N7180 Segment
X7180 N7180 N7181 Segment
X7181 N7181 N7182 Segment
X7182 N7182 N7183 Segment
X7183 N7183 N7184 Segment
X7184 N7184 N7185 Segment
X7185 N7185 N7186 Segment
X7186 N7186 N7187 Segment
X7187 N7187 N7188 Segment
X7188 N7188 N7189 Segment
X7189 N7189 N7190 Segment
X7190 N7190 N7191 Segment
X7191 N7191 N7192 Segment
X7192 N7192 N7193 Segment
X7193 N7193 N7194 Segment
X7194 N7194 N7195 Segment
X7195 N7195 N7196 Segment
X7196 N7196 N7197 Segment
X7197 N7197 N7198 Segment
X7198 N7198 N7199 Segment
X7199 N7199 N7200 Segment
X7200 N7200 N7201 Segment
X7201 N7201 N7202 Segment
X7202 N7202 N7203 Segment
X7203 N7203 N7204 Segment
X7204 N7204 N7205 Segment
X7205 N7205 N7206 Segment
X7206 N7206 N7207 Segment
X7207 N7207 N7208 Segment
X7208 N7208 N7209 Segment
X7209 N7209 N7210 Segment
X7210 N7210 N7211 Segment
X7211 N7211 N7212 Segment
X7212 N7212 N7213 Segment
X7213 N7213 N7214 Segment
X7214 N7214 N7215 Segment
X7215 N7215 N7216 Segment
X7216 N7216 N7217 Segment
X7217 N7217 N7218 Segment
X7218 N7218 N7219 Segment
X7219 N7219 N7220 Segment
X7220 N7220 N7221 Segment
X7221 N7221 N7222 Segment
X7222 N7222 N7223 Segment
X7223 N7223 N7224 Segment
X7224 N7224 N7225 Segment
X7225 N7225 N7226 Segment
X7226 N7226 N7227 Segment
X7227 N7227 N7228 Segment
X7228 N7228 N7229 Segment
X7229 N7229 N7230 Segment
X7230 N7230 N7231 Segment
X7231 N7231 N7232 Segment
X7232 N7232 N7233 Segment
X7233 N7233 N7234 Segment
X7234 N7234 N7235 Segment
X7235 N7235 N7236 Segment
X7236 N7236 N7237 Segment
X7237 N7237 N7238 Segment
X7238 N7238 N7239 Segment
X7239 N7239 N7240 Segment
X7240 N7240 N7241 Segment
X7241 N7241 N7242 Segment
X7242 N7242 N7243 Segment
X7243 N7243 N7244 Segment
X7244 N7244 N7245 Segment
X7245 N7245 N7246 Segment
X7246 N7246 N7247 Segment
X7247 N7247 N7248 Segment
X7248 N7248 N7249 Segment
X7249 N7249 N7250 Segment
X7250 N7250 N7251 Segment
X7251 N7251 N7252 Segment
X7252 N7252 N7253 Segment
X7253 N7253 N7254 Segment
X7254 N7254 N7255 Segment
X7255 N7255 N7256 Segment
X7256 N7256 N7257 Segment
X7257 N7257 N7258 Segment
X7258 N7258 N7259 Segment
X7259 N7259 N7260 Segment
X7260 N7260 N7261 Segment
X7261 N7261 N7262 Segment
X7262 N7262 N7263 Segment
X7263 N7263 N7264 Segment
X7264 N7264 N7265 Segment
X7265 N7265 N7266 Segment
X7266 N7266 N7267 Segment
X7267 N7267 N7268 Segment
X7268 N7268 N7269 Segment
X7269 N7269 N7270 Segment
X7270 N7270 N7271 Segment
X7271 N7271 N7272 Segment
X7272 N7272 N7273 Segment
X7273 N7273 N7274 Segment
X7274 N7274 N7275 Segment
X7275 N7275 N7276 Segment
X7276 N7276 N7277 Segment
X7277 N7277 N7278 Segment
X7278 N7278 N7279 Segment
X7279 N7279 N7280 Segment
X7280 N7280 N7281 Segment
X7281 N7281 N7282 Segment
X7282 N7282 N7283 Segment
X7283 N7283 N7284 Segment
X7284 N7284 N7285 Segment
X7285 N7285 N7286 Segment
X7286 N7286 N7287 Segment
X7287 N7287 N7288 Segment
X7288 N7288 N7289 Segment
X7289 N7289 N7290 Segment
X7290 N7290 N7291 Segment
X7291 N7291 N7292 Segment
X7292 N7292 N7293 Segment
X7293 N7293 N7294 Segment
X7294 N7294 N7295 Segment
X7295 N7295 N7296 Segment
X7296 N7296 N7297 Segment
X7297 N7297 N7298 Segment
X7298 N7298 N7299 Segment
X7299 N7299 N7300 Segment
X7300 N7300 N7301 Segment
X7301 N7301 N7302 Segment
X7302 N7302 N7303 Segment
X7303 N7303 N7304 Segment
X7304 N7304 N7305 Segment
X7305 N7305 N7306 Segment
X7306 N7306 N7307 Segment
X7307 N7307 N7308 Segment
X7308 N7308 N7309 Segment
X7309 N7309 N7310 Segment
X7310 N7310 N7311 Segment
X7311 N7311 N7312 Segment
X7312 N7312 N7313 Segment
X7313 N7313 N7314 Segment
X7314 N7314 N7315 Segment
X7315 N7315 N7316 Segment
X7316 N7316 N7317 Segment
X7317 N7317 N7318 Segment
X7318 N7318 N7319 Segment
X7319 N7319 N7320 Segment
X7320 N7320 N7321 Segment
X7321 N7321 N7322 Segment
X7322 N7322 N7323 Segment
X7323 N7323 N7324 Segment
X7324 N7324 N7325 Segment
X7325 N7325 N7326 Segment
X7326 N7326 N7327 Segment
X7327 N7327 N7328 Segment
X7328 N7328 N7329 Segment
X7329 N7329 N7330 Segment
X7330 N7330 N7331 Segment
X7331 N7331 N7332 Segment
X7332 N7332 N7333 Segment
X7333 N7333 N7334 Segment
X7334 N7334 N7335 Segment
X7335 N7335 N7336 Segment
X7336 N7336 N7337 Segment
X7337 N7337 N7338 Segment
X7338 N7338 N7339 Segment
X7339 N7339 N7340 Segment
X7340 N7340 N7341 Segment
X7341 N7341 N7342 Segment
X7342 N7342 N7343 Segment
X7343 N7343 N7344 Segment
X7344 N7344 N7345 Segment
X7345 N7345 N7346 Segment
X7346 N7346 N7347 Segment
X7347 N7347 N7348 Segment
X7348 N7348 N7349 Segment
X7349 N7349 N7350 Segment
X7350 N7350 N7351 Segment
X7351 N7351 N7352 Segment
X7352 N7352 N7353 Segment
X7353 N7353 N7354 Segment
X7354 N7354 N7355 Segment
X7355 N7355 N7356 Segment
X7356 N7356 N7357 Segment
X7357 N7357 N7358 Segment
X7358 N7358 N7359 Segment
X7359 N7359 N7360 Segment
X7360 N7360 N7361 Segment
X7361 N7361 N7362 Segment
X7362 N7362 N7363 Segment
X7363 N7363 N7364 Segment
X7364 N7364 N7365 Segment
X7365 N7365 N7366 Segment
X7366 N7366 N7367 Segment
X7367 N7367 N7368 Segment
X7368 N7368 N7369 Segment
X7369 N7369 N7370 Segment
X7370 N7370 N7371 Segment
X7371 N7371 N7372 Segment
X7372 N7372 N7373 Segment
X7373 N7373 N7374 Segment
X7374 N7374 N7375 Segment
X7375 N7375 N7376 Segment
X7376 N7376 N7377 Segment
X7377 N7377 N7378 Segment
X7378 N7378 N7379 Segment
X7379 N7379 N7380 Segment
X7380 N7380 N7381 Segment
X7381 N7381 N7382 Segment
X7382 N7382 N7383 Segment
X7383 N7383 N7384 Segment
X7384 N7384 N7385 Segment
X7385 N7385 N7386 Segment
X7386 N7386 N7387 Segment
X7387 N7387 N7388 Segment
X7388 N7388 N7389 Segment
X7389 N7389 N7390 Segment
X7390 N7390 N7391 Segment
X7391 N7391 N7392 Segment
X7392 N7392 N7393 Segment
X7393 N7393 N7394 Segment
X7394 N7394 N7395 Segment
X7395 N7395 N7396 Segment
X7396 N7396 N7397 Segment
X7397 N7397 N7398 Segment
X7398 N7398 N7399 Segment
X7399 N7399 N7400 Segment
X7400 N7400 N7401 Segment
X7401 N7401 N7402 Segment
X7402 N7402 N7403 Segment
X7403 N7403 N7404 Segment
X7404 N7404 N7405 Segment
X7405 N7405 N7406 Segment
X7406 N7406 N7407 Segment
X7407 N7407 N7408 Segment
X7408 N7408 N7409 Segment
X7409 N7409 N7410 Segment
X7410 N7410 N7411 Segment
X7411 N7411 N7412 Segment
X7412 N7412 N7413 Segment
X7413 N7413 N7414 Segment
X7414 N7414 N7415 Segment
X7415 N7415 N7416 Segment
X7416 N7416 N7417 Segment
X7417 N7417 N7418 Segment
X7418 N7418 N7419 Segment
X7419 N7419 N7420 Segment
X7420 N7420 N7421 Segment
X7421 N7421 N7422 Segment
X7422 N7422 N7423 Segment
X7423 N7423 N7424 Segment
X7424 N7424 N7425 Segment
X7425 N7425 N7426 Segment
X7426 N7426 N7427 Segment
X7427 N7427 N7428 Segment
X7428 N7428 N7429 Segment
X7429 N7429 N7430 Segment
X7430 N7430 N7431 Segment
X7431 N7431 N7432 Segment
X7432 N7432 N7433 Segment
X7433 N7433 N7434 Segment
X7434 N7434 N7435 Segment
X7435 N7435 N7436 Segment
X7436 N7436 N7437 Segment
X7437 N7437 N7438 Segment
X7438 N7438 N7439 Segment
X7439 N7439 N7440 Segment
X7440 N7440 N7441 Segment
X7441 N7441 N7442 Segment
X7442 N7442 N7443 Segment
X7443 N7443 N7444 Segment
X7444 N7444 N7445 Segment
X7445 N7445 N7446 Segment
X7446 N7446 N7447 Segment
X7447 N7447 N7448 Segment
X7448 N7448 N7449 Segment
X7449 N7449 N7450 Segment
X7450 N7450 N7451 Segment
X7451 N7451 N7452 Segment
X7452 N7452 N7453 Segment
X7453 N7453 N7454 Segment
X7454 N7454 N7455 Segment
X7455 N7455 N7456 Segment
X7456 N7456 N7457 Segment
X7457 N7457 N7458 Segment
X7458 N7458 N7459 Segment
X7459 N7459 N7460 Segment
X7460 N7460 N7461 Segment
X7461 N7461 N7462 Segment
X7462 N7462 N7463 Segment
X7463 N7463 N7464 Segment
X7464 N7464 N7465 Segment
X7465 N7465 N7466 Segment
X7466 N7466 N7467 Segment
X7467 N7467 N7468 Segment
X7468 N7468 N7469 Segment
X7469 N7469 N7470 Segment
X7470 N7470 N7471 Segment
X7471 N7471 N7472 Segment
X7472 N7472 N7473 Segment
X7473 N7473 N7474 Segment
X7474 N7474 N7475 Segment
X7475 N7475 N7476 Segment
X7476 N7476 N7477 Segment
X7477 N7477 N7478 Segment
X7478 N7478 N7479 Segment
X7479 N7479 N7480 Segment
X7480 N7480 N7481 Segment
X7481 N7481 N7482 Segment
X7482 N7482 N7483 Segment
X7483 N7483 N7484 Segment
X7484 N7484 N7485 Segment
X7485 N7485 N7486 Segment
X7486 N7486 N7487 Segment
X7487 N7487 N7488 Segment
X7488 N7488 N7489 Segment
X7489 N7489 N7490 Segment
X7490 N7490 N7491 Segment
X7491 N7491 N7492 Segment
X7492 N7492 N7493 Segment
X7493 N7493 N7494 Segment
X7494 N7494 N7495 Segment
X7495 N7495 N7496 Segment
X7496 N7496 N7497 Segment
X7497 N7497 N7498 Segment
X7498 N7498 N7499 Segment
X7499 N7499 N7500 Segment
X7500 N7500 N7501 Segment
X7501 N7501 N7502 Segment
X7502 N7502 N7503 Segment
X7503 N7503 N7504 Segment
X7504 N7504 N7505 Segment
X7505 N7505 N7506 Segment
X7506 N7506 N7507 Segment
X7507 N7507 N7508 Segment
X7508 N7508 N7509 Segment
X7509 N7509 N7510 Segment
X7510 N7510 N7511 Segment
X7511 N7511 N7512 Segment
X7512 N7512 N7513 Segment
X7513 N7513 N7514 Segment
X7514 N7514 N7515 Segment
X7515 N7515 N7516 Segment
X7516 N7516 N7517 Segment
X7517 N7517 N7518 Segment
X7518 N7518 N7519 Segment
X7519 N7519 N7520 Segment
X7520 N7520 N7521 Segment
X7521 N7521 N7522 Segment
X7522 N7522 N7523 Segment
X7523 N7523 N7524 Segment
X7524 N7524 N7525 Segment
X7525 N7525 N7526 Segment
X7526 N7526 N7527 Segment
X7527 N7527 N7528 Segment
X7528 N7528 N7529 Segment
X7529 N7529 N7530 Segment
X7530 N7530 N7531 Segment
X7531 N7531 N7532 Segment
X7532 N7532 N7533 Segment
X7533 N7533 N7534 Segment
X7534 N7534 N7535 Segment
X7535 N7535 N7536 Segment
X7536 N7536 N7537 Segment
X7537 N7537 N7538 Segment
X7538 N7538 N7539 Segment
X7539 N7539 N7540 Segment
X7540 N7540 N7541 Segment
X7541 N7541 N7542 Segment
X7542 N7542 N7543 Segment
X7543 N7543 N7544 Segment
X7544 N7544 N7545 Segment
X7545 N7545 N7546 Segment
X7546 N7546 N7547 Segment
X7547 N7547 N7548 Segment
X7548 N7548 N7549 Segment
X7549 N7549 N7550 Segment
X7550 N7550 N7551 Segment
X7551 N7551 N7552 Segment
X7552 N7552 N7553 Segment
X7553 N7553 N7554 Segment
X7554 N7554 N7555 Segment
X7555 N7555 N7556 Segment
X7556 N7556 N7557 Segment
X7557 N7557 N7558 Segment
X7558 N7558 N7559 Segment
X7559 N7559 N7560 Segment
X7560 N7560 N7561 Segment
X7561 N7561 N7562 Segment
X7562 N7562 N7563 Segment
X7563 N7563 N7564 Segment
X7564 N7564 N7565 Segment
X7565 N7565 N7566 Segment
X7566 N7566 N7567 Segment
X7567 N7567 N7568 Segment
X7568 N7568 N7569 Segment
X7569 N7569 N7570 Segment
X7570 N7570 N7571 Segment
X7571 N7571 N7572 Segment
X7572 N7572 N7573 Segment
X7573 N7573 N7574 Segment
X7574 N7574 N7575 Segment
X7575 N7575 N7576 Segment
X7576 N7576 N7577 Segment
X7577 N7577 N7578 Segment
X7578 N7578 N7579 Segment
X7579 N7579 N7580 Segment
X7580 N7580 N7581 Segment
X7581 N7581 N7582 Segment
X7582 N7582 N7583 Segment
X7583 N7583 N7584 Segment
X7584 N7584 N7585 Segment
X7585 N7585 N7586 Segment
X7586 N7586 N7587 Segment
X7587 N7587 N7588 Segment
X7588 N7588 N7589 Segment
X7589 N7589 N7590 Segment
X7590 N7590 N7591 Segment
X7591 N7591 N7592 Segment
X7592 N7592 N7593 Segment
X7593 N7593 N7594 Segment
X7594 N7594 N7595 Segment
X7595 N7595 N7596 Segment
X7596 N7596 N7597 Segment
X7597 N7597 N7598 Segment
X7598 N7598 N7599 Segment
X7599 N7599 N7600 Segment
X7600 N7600 N7601 Segment
X7601 N7601 N7602 Segment
X7602 N7602 N7603 Segment
X7603 N7603 N7604 Segment
X7604 N7604 N7605 Segment
X7605 N7605 N7606 Segment
X7606 N7606 N7607 Segment
X7607 N7607 N7608 Segment
X7608 N7608 N7609 Segment
X7609 N7609 N7610 Segment
X7610 N7610 N7611 Segment
X7611 N7611 N7612 Segment
X7612 N7612 N7613 Segment
X7613 N7613 N7614 Segment
X7614 N7614 N7615 Segment
X7615 N7615 N7616 Segment
X7616 N7616 N7617 Segment
X7617 N7617 N7618 Segment
X7618 N7618 N7619 Segment
X7619 N7619 N7620 Segment
X7620 N7620 N7621 Segment
X7621 N7621 N7622 Segment
X7622 N7622 N7623 Segment
X7623 N7623 N7624 Segment
X7624 N7624 N7625 Segment
X7625 N7625 N7626 Segment
X7626 N7626 N7627 Segment
X7627 N7627 N7628 Segment
X7628 N7628 N7629 Segment
X7629 N7629 N7630 Segment
X7630 N7630 N7631 Segment
X7631 N7631 N7632 Segment
X7632 N7632 N7633 Segment
X7633 N7633 N7634 Segment
X7634 N7634 N7635 Segment
X7635 N7635 N7636 Segment
X7636 N7636 N7637 Segment
X7637 N7637 N7638 Segment
X7638 N7638 N7639 Segment
X7639 N7639 N7640 Segment
X7640 N7640 N7641 Segment
X7641 N7641 N7642 Segment
X7642 N7642 N7643 Segment
X7643 N7643 N7644 Segment
X7644 N7644 N7645 Segment
X7645 N7645 N7646 Segment
X7646 N7646 N7647 Segment
X7647 N7647 N7648 Segment
X7648 N7648 N7649 Segment
X7649 N7649 N7650 Segment
X7650 N7650 N7651 Segment
X7651 N7651 N7652 Segment
X7652 N7652 N7653 Segment
X7653 N7653 N7654 Segment
X7654 N7654 N7655 Segment
X7655 N7655 N7656 Segment
X7656 N7656 N7657 Segment
X7657 N7657 N7658 Segment
X7658 N7658 N7659 Segment
X7659 N7659 N7660 Segment
X7660 N7660 N7661 Segment
X7661 N7661 N7662 Segment
X7662 N7662 N7663 Segment
X7663 N7663 N7664 Segment
X7664 N7664 N7665 Segment
X7665 N7665 N7666 Segment
X7666 N7666 N7667 Segment
X7667 N7667 N7668 Segment
X7668 N7668 N7669 Segment
X7669 N7669 N7670 Segment
X7670 N7670 N7671 Segment
X7671 N7671 N7672 Segment
X7672 N7672 N7673 Segment
X7673 N7673 N7674 Segment
X7674 N7674 N7675 Segment
X7675 N7675 N7676 Segment
X7676 N7676 N7677 Segment
X7677 N7677 N7678 Segment
X7678 N7678 N7679 Segment
X7679 N7679 N7680 Segment
X7680 N7680 N7681 Segment
X7681 N7681 N7682 Segment
X7682 N7682 N7683 Segment
X7683 N7683 N7684 Segment
X7684 N7684 N7685 Segment
X7685 N7685 N7686 Segment
X7686 N7686 N7687 Segment
X7687 N7687 N7688 Segment
X7688 N7688 N7689 Segment
X7689 N7689 N7690 Segment
X7690 N7690 N7691 Segment
X7691 N7691 N7692 Segment
X7692 N7692 N7693 Segment
X7693 N7693 N7694 Segment
X7694 N7694 N7695 Segment
X7695 N7695 N7696 Segment
X7696 N7696 N7697 Segment
X7697 N7697 N7698 Segment
X7698 N7698 N7699 Segment
X7699 N7699 N7700 Segment
X7700 N7700 N7701 Segment
X7701 N7701 N7702 Segment
X7702 N7702 N7703 Segment
X7703 N7703 N7704 Segment
X7704 N7704 N7705 Segment
X7705 N7705 N7706 Segment
X7706 N7706 N7707 Segment
X7707 N7707 N7708 Segment
X7708 N7708 N7709 Segment
X7709 N7709 N7710 Segment
X7710 N7710 N7711 Segment
X7711 N7711 N7712 Segment
X7712 N7712 N7713 Segment
X7713 N7713 N7714 Segment
X7714 N7714 N7715 Segment
X7715 N7715 N7716 Segment
X7716 N7716 N7717 Segment
X7717 N7717 N7718 Segment
X7718 N7718 N7719 Segment
X7719 N7719 N7720 Segment
X7720 N7720 N7721 Segment
X7721 N7721 N7722 Segment
X7722 N7722 N7723 Segment
X7723 N7723 N7724 Segment
X7724 N7724 N7725 Segment
X7725 N7725 N7726 Segment
X7726 N7726 N7727 Segment
X7727 N7727 N7728 Segment
X7728 N7728 N7729 Segment
X7729 N7729 N7730 Segment
X7730 N7730 N7731 Segment
X7731 N7731 N7732 Segment
X7732 N7732 N7733 Segment
X7733 N7733 N7734 Segment
X7734 N7734 N7735 Segment
X7735 N7735 N7736 Segment
X7736 N7736 N7737 Segment
X7737 N7737 N7738 Segment
X7738 N7738 N7739 Segment
X7739 N7739 N7740 Segment
X7740 N7740 N7741 Segment
X7741 N7741 N7742 Segment
X7742 N7742 N7743 Segment
X7743 N7743 N7744 Segment
X7744 N7744 N7745 Segment
X7745 N7745 N7746 Segment
X7746 N7746 N7747 Segment
X7747 N7747 N7748 Segment
X7748 N7748 N7749 Segment
X7749 N7749 N7750 Segment
X7750 N7750 N7751 Segment
X7751 N7751 N7752 Segment
X7752 N7752 N7753 Segment
X7753 N7753 N7754 Segment
X7754 N7754 N7755 Segment
X7755 N7755 N7756 Segment
X7756 N7756 N7757 Segment
X7757 N7757 N7758 Segment
X7758 N7758 N7759 Segment
X7759 N7759 N7760 Segment
X7760 N7760 N7761 Segment
X7761 N7761 N7762 Segment
X7762 N7762 N7763 Segment
X7763 N7763 N7764 Segment
X7764 N7764 N7765 Segment
X7765 N7765 N7766 Segment
X7766 N7766 N7767 Segment
X7767 N7767 N7768 Segment
X7768 N7768 N7769 Segment
X7769 N7769 N7770 Segment
X7770 N7770 N7771 Segment
X7771 N7771 N7772 Segment
X7772 N7772 N7773 Segment
X7773 N7773 N7774 Segment
X7774 N7774 N7775 Segment
X7775 N7775 N7776 Segment
X7776 N7776 N7777 Segment
X7777 N7777 N7778 Segment
X7778 N7778 N7779 Segment
X7779 N7779 N7780 Segment
X7780 N7780 N7781 Segment
X7781 N7781 N7782 Segment
X7782 N7782 N7783 Segment
X7783 N7783 N7784 Segment
X7784 N7784 N7785 Segment
X7785 N7785 N7786 Segment
X7786 N7786 N7787 Segment
X7787 N7787 N7788 Segment
X7788 N7788 N7789 Segment
X7789 N7789 N7790 Segment
X7790 N7790 N7791 Segment
X7791 N7791 N7792 Segment
X7792 N7792 N7793 Segment
X7793 N7793 N7794 Segment
X7794 N7794 N7795 Segment
X7795 N7795 N7796 Segment
X7796 N7796 N7797 Segment
X7797 N7797 N7798 Segment
X7798 N7798 N7799 Segment
X7799 N7799 N7800 Segment
X7800 N7800 N7801 Segment
X7801 N7801 N7802 Segment
X7802 N7802 N7803 Segment
X7803 N7803 N7804 Segment
X7804 N7804 N7805 Segment
X7805 N7805 N7806 Segment
X7806 N7806 N7807 Segment
X7807 N7807 N7808 Segment
X7808 N7808 N7809 Segment
X7809 N7809 N7810 Segment
X7810 N7810 N7811 Segment
X7811 N7811 N7812 Segment
X7812 N7812 N7813 Segment
X7813 N7813 N7814 Segment
X7814 N7814 N7815 Segment
X7815 N7815 N7816 Segment
X7816 N7816 N7817 Segment
X7817 N7817 N7818 Segment
X7818 N7818 N7819 Segment
X7819 N7819 N7820 Segment
X7820 N7820 N7821 Segment
X7821 N7821 N7822 Segment
X7822 N7822 N7823 Segment
X7823 N7823 N7824 Segment
X7824 N7824 N7825 Segment
X7825 N7825 N7826 Segment
X7826 N7826 N7827 Segment
X7827 N7827 N7828 Segment
X7828 N7828 N7829 Segment
X7829 N7829 N7830 Segment
X7830 N7830 N7831 Segment
X7831 N7831 N7832 Segment
X7832 N7832 N7833 Segment
X7833 N7833 N7834 Segment
X7834 N7834 N7835 Segment
X7835 N7835 N7836 Segment
X7836 N7836 N7837 Segment
X7837 N7837 N7838 Segment
X7838 N7838 N7839 Segment
X7839 N7839 N7840 Segment
X7840 N7840 N7841 Segment
X7841 N7841 N7842 Segment
X7842 N7842 N7843 Segment
X7843 N7843 N7844 Segment
X7844 N7844 N7845 Segment
X7845 N7845 N7846 Segment
X7846 N7846 N7847 Segment
X7847 N7847 N7848 Segment
X7848 N7848 N7849 Segment
X7849 N7849 N7850 Segment
X7850 N7850 N7851 Segment
X7851 N7851 N7852 Segment
X7852 N7852 N7853 Segment
X7853 N7853 N7854 Segment
X7854 N7854 N7855 Segment
X7855 N7855 N7856 Segment
X7856 N7856 N7857 Segment
X7857 N7857 N7858 Segment
X7858 N7858 N7859 Segment
X7859 N7859 N7860 Segment
X7860 N7860 N7861 Segment
X7861 N7861 N7862 Segment
X7862 N7862 N7863 Segment
X7863 N7863 N7864 Segment
X7864 N7864 N7865 Segment
X7865 N7865 N7866 Segment
X7866 N7866 N7867 Segment
X7867 N7867 N7868 Segment
X7868 N7868 N7869 Segment
X7869 N7869 N7870 Segment
X7870 N7870 N7871 Segment
X7871 N7871 N7872 Segment
X7872 N7872 N7873 Segment
X7873 N7873 N7874 Segment
X7874 N7874 N7875 Segment
X7875 N7875 N7876 Segment
X7876 N7876 N7877 Segment
X7877 N7877 N7878 Segment
X7878 N7878 N7879 Segment
X7879 N7879 N7880 Segment
X7880 N7880 N7881 Segment
X7881 N7881 N7882 Segment
X7882 N7882 N7883 Segment
X7883 N7883 N7884 Segment
X7884 N7884 N7885 Segment
X7885 N7885 N7886 Segment
X7886 N7886 N7887 Segment
X7887 N7887 N7888 Segment
X7888 N7888 N7889 Segment
X7889 N7889 N7890 Segment
X7890 N7890 N7891 Segment
X7891 N7891 N7892 Segment
X7892 N7892 N7893 Segment
X7893 N7893 N7894 Segment
X7894 N7894 N7895 Segment
X7895 N7895 N7896 Segment
X7896 N7896 N7897 Segment
X7897 N7897 N7898 Segment
X7898 N7898 N7899 Segment
X7899 N7899 N7900 Segment
X7900 N7900 N7901 Segment
X7901 N7901 N7902 Segment
X7902 N7902 N7903 Segment
X7903 N7903 N7904 Segment
X7904 N7904 N7905 Segment
X7905 N7905 N7906 Segment
X7906 N7906 N7907 Segment
X7907 N7907 N7908 Segment
X7908 N7908 N7909 Segment
X7909 N7909 N7910 Segment
X7910 N7910 N7911 Segment
X7911 N7911 N7912 Segment
X7912 N7912 N7913 Segment
X7913 N7913 N7914 Segment
X7914 N7914 N7915 Segment
X7915 N7915 N7916 Segment
X7916 N7916 N7917 Segment
X7917 N7917 N7918 Segment
X7918 N7918 N7919 Segment
X7919 N7919 N7920 Segment
X7920 N7920 N7921 Segment
X7921 N7921 N7922 Segment
X7922 N7922 N7923 Segment
X7923 N7923 N7924 Segment
X7924 N7924 N7925 Segment
X7925 N7925 N7926 Segment
X7926 N7926 N7927 Segment
X7927 N7927 N7928 Segment
X7928 N7928 N7929 Segment
X7929 N7929 N7930 Segment
X7930 N7930 N7931 Segment
X7931 N7931 N7932 Segment
X7932 N7932 N7933 Segment
X7933 N7933 N7934 Segment
X7934 N7934 N7935 Segment
X7935 N7935 N7936 Segment
X7936 N7936 N7937 Segment
X7937 N7937 N7938 Segment
X7938 N7938 N7939 Segment
X7939 N7939 N7940 Segment
X7940 N7940 N7941 Segment
X7941 N7941 N7942 Segment
X7942 N7942 N7943 Segment
X7943 N7943 N7944 Segment
X7944 N7944 N7945 Segment
X7945 N7945 N7946 Segment
X7946 N7946 N7947 Segment
X7947 N7947 N7948 Segment
X7948 N7948 N7949 Segment
X7949 N7949 N7950 Segment
X7950 N7950 N7951 Segment
X7951 N7951 N7952 Segment
X7952 N7952 N7953 Segment
X7953 N7953 N7954 Segment
X7954 N7954 N7955 Segment
X7955 N7955 N7956 Segment
X7956 N7956 N7957 Segment
X7957 N7957 N7958 Segment
X7958 N7958 N7959 Segment
X7959 N7959 N7960 Segment
X7960 N7960 N7961 Segment
X7961 N7961 N7962 Segment
X7962 N7962 N7963 Segment
X7963 N7963 N7964 Segment
X7964 N7964 N7965 Segment
X7965 N7965 N7966 Segment
X7966 N7966 N7967 Segment
X7967 N7967 N7968 Segment
X7968 N7968 N7969 Segment
X7969 N7969 N7970 Segment
X7970 N7970 N7971 Segment
X7971 N7971 N7972 Segment
X7972 N7972 N7973 Segment
X7973 N7973 N7974 Segment
X7974 N7974 N7975 Segment
X7975 N7975 N7976 Segment
X7976 N7976 N7977 Segment
X7977 N7977 N7978 Segment
X7978 N7978 N7979 Segment
X7979 N7979 N7980 Segment
X7980 N7980 N7981 Segment
X7981 N7981 N7982 Segment
X7982 N7982 N7983 Segment
X7983 N7983 N7984 Segment
X7984 N7984 N7985 Segment
X7985 N7985 N7986 Segment
X7986 N7986 N7987 Segment
X7987 N7987 N7988 Segment
X7988 N7988 N7989 Segment
X7989 N7989 N7990 Segment
X7990 N7990 N7991 Segment
X7991 N7991 N7992 Segment
X7992 N7992 N7993 Segment
X7993 N7993 N7994 Segment
X7994 N7994 N7995 Segment
X7995 N7995 N7996 Segment
X7996 N7996 N7997 Segment
X7997 N7997 N7998 Segment
X7998 N7998 N7999 Segment
X7999 N7999 N8000 Segment
X8000 N8000 N8001 Segment
X8001 N8001 N8002 Segment
X8002 N8002 N8003 Segment
X8003 N8003 N8004 Segment
X8004 N8004 N8005 Segment
X8005 N8005 N8006 Segment
X8006 N8006 N8007 Segment
X8007 N8007 N8008 Segment
X8008 N8008 N8009 Segment
X8009 N8009 N8010 Segment
X8010 N8010 N8011 Segment
X8011 N8011 N8012 Segment
X8012 N8012 N8013 Segment
X8013 N8013 N8014 Segment
X8014 N8014 N8015 Segment
X8015 N8015 N8016 Segment
X8016 N8016 N8017 Segment
X8017 N8017 N8018 Segment
X8018 N8018 N8019 Segment
X8019 N8019 N8020 Segment
X8020 N8020 N8021 Segment
X8021 N8021 N8022 Segment
X8022 N8022 N8023 Segment
X8023 N8023 N8024 Segment
X8024 N8024 N8025 Segment
X8025 N8025 N8026 Segment
X8026 N8026 N8027 Segment
X8027 N8027 N8028 Segment
X8028 N8028 N8029 Segment
X8029 N8029 N8030 Segment
X8030 N8030 N8031 Segment
X8031 N8031 N8032 Segment
X8032 N8032 N8033 Segment
X8033 N8033 N8034 Segment
X8034 N8034 N8035 Segment
X8035 N8035 N8036 Segment
X8036 N8036 N8037 Segment
X8037 N8037 N8038 Segment
X8038 N8038 N8039 Segment
X8039 N8039 N8040 Segment
X8040 N8040 N8041 Segment
X8041 N8041 N8042 Segment
X8042 N8042 N8043 Segment
X8043 N8043 N8044 Segment
X8044 N8044 N8045 Segment
X8045 N8045 N8046 Segment
X8046 N8046 N8047 Segment
X8047 N8047 N8048 Segment
X8048 N8048 N8049 Segment
X8049 N8049 N8050 Segment
X8050 N8050 N8051 Segment
X8051 N8051 N8052 Segment
X8052 N8052 N8053 Segment
X8053 N8053 N8054 Segment
X8054 N8054 N8055 Segment
X8055 N8055 N8056 Segment
X8056 N8056 N8057 Segment
X8057 N8057 N8058 Segment
X8058 N8058 N8059 Segment
X8059 N8059 N8060 Segment
X8060 N8060 N8061 Segment
X8061 N8061 N8062 Segment
X8062 N8062 N8063 Segment
X8063 N8063 N8064 Segment
X8064 N8064 N8065 Segment
X8065 N8065 N8066 Segment
X8066 N8066 N8067 Segment
X8067 N8067 N8068 Segment
X8068 N8068 N8069 Segment
X8069 N8069 N8070 Segment
X8070 N8070 N8071 Segment
X8071 N8071 N8072 Segment
X8072 N8072 N8073 Segment
X8073 N8073 N8074 Segment
X8074 N8074 N8075 Segment
X8075 N8075 N8076 Segment
X8076 N8076 N8077 Segment
X8077 N8077 N8078 Segment
X8078 N8078 N8079 Segment
X8079 N8079 N8080 Segment
X8080 N8080 N8081 Segment
X8081 N8081 N8082 Segment
X8082 N8082 N8083 Segment
X8083 N8083 N8084 Segment
X8084 N8084 N8085 Segment
X8085 N8085 N8086 Segment
X8086 N8086 N8087 Segment
X8087 N8087 N8088 Segment
X8088 N8088 N8089 Segment
X8089 N8089 N8090 Segment
X8090 N8090 N8091 Segment
X8091 N8091 N8092 Segment
X8092 N8092 N8093 Segment
X8093 N8093 N8094 Segment
X8094 N8094 N8095 Segment
X8095 N8095 N8096 Segment
X8096 N8096 N8097 Segment
X8097 N8097 N8098 Segment
X8098 N8098 N8099 Segment
X8099 N8099 N8100 Segment
X8100 N8100 N8101 Segment
X8101 N8101 N8102 Segment
X8102 N8102 N8103 Segment
X8103 N8103 N8104 Segment
X8104 N8104 N8105 Segment
X8105 N8105 N8106 Segment
X8106 N8106 N8107 Segment
X8107 N8107 N8108 Segment
X8108 N8108 N8109 Segment
X8109 N8109 N8110 Segment
X8110 N8110 N8111 Segment
X8111 N8111 N8112 Segment
X8112 N8112 N8113 Segment
X8113 N8113 N8114 Segment
X8114 N8114 N8115 Segment
X8115 N8115 N8116 Segment
X8116 N8116 N8117 Segment
X8117 N8117 N8118 Segment
X8118 N8118 N8119 Segment
X8119 N8119 N8120 Segment
X8120 N8120 N8121 Segment
X8121 N8121 N8122 Segment
X8122 N8122 N8123 Segment
X8123 N8123 N8124 Segment
X8124 N8124 N8125 Segment
X8125 N8125 N8126 Segment
X8126 N8126 N8127 Segment
X8127 N8127 N8128 Segment
X8128 N8128 N8129 Segment
X8129 N8129 N8130 Segment
X8130 N8130 N8131 Segment
X8131 N8131 N8132 Segment
X8132 N8132 N8133 Segment
X8133 N8133 N8134 Segment
X8134 N8134 N8135 Segment
X8135 N8135 N8136 Segment
X8136 N8136 N8137 Segment
X8137 N8137 N8138 Segment
X8138 N8138 N8139 Segment
X8139 N8139 N8140 Segment
X8140 N8140 N8141 Segment
X8141 N8141 N8142 Segment
X8142 N8142 N8143 Segment
X8143 N8143 N8144 Segment
X8144 N8144 N8145 Segment
X8145 N8145 N8146 Segment
X8146 N8146 N8147 Segment
X8147 N8147 N8148 Segment
X8148 N8148 N8149 Segment
X8149 N8149 N8150 Segment
X8150 N8150 N8151 Segment
X8151 N8151 N8152 Segment
X8152 N8152 N8153 Segment
X8153 N8153 N8154 Segment
X8154 N8154 N8155 Segment
X8155 N8155 N8156 Segment
X8156 N8156 N8157 Segment
X8157 N8157 N8158 Segment
X8158 N8158 N8159 Segment
X8159 N8159 N8160 Segment
X8160 N8160 N8161 Segment
X8161 N8161 N8162 Segment
X8162 N8162 N8163 Segment
X8163 N8163 N8164 Segment
X8164 N8164 N8165 Segment
X8165 N8165 N8166 Segment
X8166 N8166 N8167 Segment
X8167 N8167 N8168 Segment
X8168 N8168 N8169 Segment
X8169 N8169 N8170 Segment
X8170 N8170 N8171 Segment
X8171 N8171 N8172 Segment
X8172 N8172 N8173 Segment
X8173 N8173 N8174 Segment
X8174 N8174 N8175 Segment
X8175 N8175 N8176 Segment
X8176 N8176 N8177 Segment
X8177 N8177 N8178 Segment
X8178 N8178 N8179 Segment
X8179 N8179 N8180 Segment
X8180 N8180 N8181 Segment
X8181 N8181 N8182 Segment
X8182 N8182 N8183 Segment
X8183 N8183 N8184 Segment
X8184 N8184 N8185 Segment
X8185 N8185 N8186 Segment
X8186 N8186 N8187 Segment
X8187 N8187 N8188 Segment
X8188 N8188 N8189 Segment
X8189 N8189 N8190 Segment
X8190 N8190 N8191 Segment
X8191 N8191 N8192 Segment
X8192 N8192 N8193 Segment
X8193 N8193 N8194 Segment
X8194 N8194 N8195 Segment
X8195 N8195 N8196 Segment
X8196 N8196 N8197 Segment
X8197 N8197 N8198 Segment
X8198 N8198 N8199 Segment
X8199 N8199 N8200 Segment
X8200 N8200 N8201 Segment
X8201 N8201 N8202 Segment
X8202 N8202 N8203 Segment
X8203 N8203 N8204 Segment
X8204 N8204 N8205 Segment
X8205 N8205 N8206 Segment
X8206 N8206 N8207 Segment
X8207 N8207 N8208 Segment
X8208 N8208 N8209 Segment
X8209 N8209 N8210 Segment
X8210 N8210 N8211 Segment
X8211 N8211 N8212 Segment
X8212 N8212 N8213 Segment
X8213 N8213 N8214 Segment
X8214 N8214 N8215 Segment
X8215 N8215 N8216 Segment
X8216 N8216 N8217 Segment
X8217 N8217 N8218 Segment
X8218 N8218 N8219 Segment
X8219 N8219 N8220 Segment
X8220 N8220 N8221 Segment
X8221 N8221 N8222 Segment
X8222 N8222 N8223 Segment
X8223 N8223 N8224 Segment
X8224 N8224 N8225 Segment
X8225 N8225 N8226 Segment
X8226 N8226 N8227 Segment
X8227 N8227 N8228 Segment
X8228 N8228 N8229 Segment
X8229 N8229 N8230 Segment
X8230 N8230 N8231 Segment
X8231 N8231 N8232 Segment
X8232 N8232 N8233 Segment
X8233 N8233 N8234 Segment
X8234 N8234 N8235 Segment
X8235 N8235 N8236 Segment
X8236 N8236 N8237 Segment
X8237 N8237 N8238 Segment
X8238 N8238 N8239 Segment
X8239 N8239 N8240 Segment
X8240 N8240 N8241 Segment
X8241 N8241 N8242 Segment
X8242 N8242 N8243 Segment
X8243 N8243 N8244 Segment
X8244 N8244 N8245 Segment
X8245 N8245 N8246 Segment
X8246 N8246 N8247 Segment
X8247 N8247 N8248 Segment
X8248 N8248 N8249 Segment
X8249 N8249 N8250 Segment
X8250 N8250 N8251 Segment
X8251 N8251 N8252 Segment
X8252 N8252 N8253 Segment
X8253 N8253 N8254 Segment
X8254 N8254 N8255 Segment
X8255 N8255 N8256 Segment
X8256 N8256 N8257 Segment
X8257 N8257 N8258 Segment
X8258 N8258 N8259 Segment
X8259 N8259 N8260 Segment
X8260 N8260 N8261 Segment
X8261 N8261 N8262 Segment
X8262 N8262 N8263 Segment
X8263 N8263 N8264 Segment
X8264 N8264 N8265 Segment
X8265 N8265 N8266 Segment
X8266 N8266 N8267 Segment
X8267 N8267 N8268 Segment
X8268 N8268 N8269 Segment
X8269 N8269 N8270 Segment
X8270 N8270 N8271 Segment
X8271 N8271 N8272 Segment
X8272 N8272 N8273 Segment
X8273 N8273 N8274 Segment
X8274 N8274 N8275 Segment
X8275 N8275 N8276 Segment
X8276 N8276 N8277 Segment
X8277 N8277 N8278 Segment
X8278 N8278 N8279 Segment
X8279 N8279 N8280 Segment
X8280 N8280 N8281 Segment
X8281 N8281 N8282 Segment
X8282 N8282 N8283 Segment
X8283 N8283 N8284 Segment
X8284 N8284 N8285 Segment
X8285 N8285 N8286 Segment
X8286 N8286 N8287 Segment
X8287 N8287 N8288 Segment
X8288 N8288 N8289 Segment
X8289 N8289 N8290 Segment
X8290 N8290 N8291 Segment
X8291 N8291 N8292 Segment
X8292 N8292 N8293 Segment
X8293 N8293 N8294 Segment
X8294 N8294 N8295 Segment
X8295 N8295 N8296 Segment
X8296 N8296 N8297 Segment
X8297 N8297 N8298 Segment
X8298 N8298 N8299 Segment
X8299 N8299 N8300 Segment
X8300 N8300 N8301 Segment
X8301 N8301 N8302 Segment
X8302 N8302 N8303 Segment
X8303 N8303 N8304 Segment
X8304 N8304 N8305 Segment
X8305 N8305 N8306 Segment
X8306 N8306 N8307 Segment
X8307 N8307 N8308 Segment
X8308 N8308 N8309 Segment
X8309 N8309 N8310 Segment
X8310 N8310 N8311 Segment
X8311 N8311 N8312 Segment
X8312 N8312 N8313 Segment
X8313 N8313 N8314 Segment
X8314 N8314 N8315 Segment
X8315 N8315 N8316 Segment
X8316 N8316 N8317 Segment
X8317 N8317 N8318 Segment
X8318 N8318 N8319 Segment
X8319 N8319 N8320 Segment
X8320 N8320 N8321 Segment
X8321 N8321 N8322 Segment
X8322 N8322 N8323 Segment
X8323 N8323 N8324 Segment
X8324 N8324 N8325 Segment
X8325 N8325 N8326 Segment
X8326 N8326 N8327 Segment
X8327 N8327 N8328 Segment
X8328 N8328 N8329 Segment
X8329 N8329 N8330 Segment
X8330 N8330 N8331 Segment
X8331 N8331 N8332 Segment
X8332 N8332 N8333 Segment
X8333 N8333 N8334 Segment
X8334 N8334 N8335 Segment
X8335 N8335 N8336 Segment
X8336 N8336 N8337 Segment
X8337 N8337 N8338 Segment
X8338 N8338 N8339 Segment
X8339 N8339 N8340 Segment
X8340 N8340 N8341 Segment
X8341 N8341 N8342 Segment
X8342 N8342 N8343 Segment
X8343 N8343 N8344 Segment
X8344 N8344 N8345 Segment
X8345 N8345 N8346 Segment
X8346 N8346 N8347 Segment
X8347 N8347 N8348 Segment
X8348 N8348 N8349 Segment
X8349 N8349 N8350 Segment
X8350 N8350 N8351 Segment
X8351 N8351 N8352 Segment
X8352 N8352 N8353 Segment
X8353 N8353 N8354 Segment
X8354 N8354 N8355 Segment
X8355 N8355 N8356 Segment
X8356 N8356 N8357 Segment
X8357 N8357 N8358 Segment
X8358 N8358 N8359 Segment
X8359 N8359 N8360 Segment
X8360 N8360 N8361 Segment
X8361 N8361 N8362 Segment
X8362 N8362 N8363 Segment
X8363 N8363 N8364 Segment
X8364 N8364 N8365 Segment
X8365 N8365 N8366 Segment
X8366 N8366 N8367 Segment
X8367 N8367 N8368 Segment
X8368 N8368 N8369 Segment
X8369 N8369 N8370 Segment
X8370 N8370 N8371 Segment
X8371 N8371 N8372 Segment
X8372 N8372 N8373 Segment
X8373 N8373 N8374 Segment
X8374 N8374 N8375 Segment
X8375 N8375 N8376 Segment
X8376 N8376 N8377 Segment
X8377 N8377 N8378 Segment
X8378 N8378 N8379 Segment
X8379 N8379 N8380 Segment
X8380 N8380 N8381 Segment
X8381 N8381 N8382 Segment
X8382 N8382 N8383 Segment
X8383 N8383 N8384 Segment
X8384 N8384 N8385 Segment
X8385 N8385 N8386 Segment
X8386 N8386 N8387 Segment
X8387 N8387 N8388 Segment
X8388 N8388 N8389 Segment
X8389 N8389 N8390 Segment
X8390 N8390 N8391 Segment
X8391 N8391 N8392 Segment
X8392 N8392 N8393 Segment
X8393 N8393 N8394 Segment
X8394 N8394 N8395 Segment
X8395 N8395 N8396 Segment
X8396 N8396 N8397 Segment
X8397 N8397 N8398 Segment
X8398 N8398 N8399 Segment
X8399 N8399 N8400 Segment
X8400 N8400 N8401 Segment
X8401 N8401 N8402 Segment
X8402 N8402 N8403 Segment
X8403 N8403 N8404 Segment
X8404 N8404 N8405 Segment
X8405 N8405 N8406 Segment
X8406 N8406 N8407 Segment
X8407 N8407 N8408 Segment
X8408 N8408 N8409 Segment
X8409 N8409 N8410 Segment
X8410 N8410 N8411 Segment
X8411 N8411 N8412 Segment
X8412 N8412 N8413 Segment
X8413 N8413 N8414 Segment
X8414 N8414 N8415 Segment
X8415 N8415 N8416 Segment
X8416 N8416 N8417 Segment
X8417 N8417 N8418 Segment
X8418 N8418 N8419 Segment
X8419 N8419 N8420 Segment
X8420 N8420 N8421 Segment
X8421 N8421 N8422 Segment
X8422 N8422 N8423 Segment
X8423 N8423 N8424 Segment
X8424 N8424 N8425 Segment
X8425 N8425 N8426 Segment
X8426 N8426 N8427 Segment
X8427 N8427 N8428 Segment
X8428 N8428 N8429 Segment
X8429 N8429 N8430 Segment
X8430 N8430 N8431 Segment
X8431 N8431 N8432 Segment
X8432 N8432 N8433 Segment
X8433 N8433 N8434 Segment
X8434 N8434 N8435 Segment
X8435 N8435 N8436 Segment
X8436 N8436 N8437 Segment
X8437 N8437 N8438 Segment
X8438 N8438 N8439 Segment
X8439 N8439 N8440 Segment
X8440 N8440 N8441 Segment
X8441 N8441 N8442 Segment
X8442 N8442 N8443 Segment
X8443 N8443 N8444 Segment
X8444 N8444 N8445 Segment
X8445 N8445 N8446 Segment
X8446 N8446 N8447 Segment
X8447 N8447 N8448 Segment
X8448 N8448 N8449 Segment
X8449 N8449 N8450 Segment
X8450 N8450 N8451 Segment
X8451 N8451 N8452 Segment
X8452 N8452 N8453 Segment
X8453 N8453 N8454 Segment
X8454 N8454 N8455 Segment
X8455 N8455 N8456 Segment
X8456 N8456 N8457 Segment
X8457 N8457 N8458 Segment
X8458 N8458 N8459 Segment
X8459 N8459 N8460 Segment
X8460 N8460 N8461 Segment
X8461 N8461 N8462 Segment
X8462 N8462 N8463 Segment
X8463 N8463 N8464 Segment
X8464 N8464 N8465 Segment
X8465 N8465 N8466 Segment
X8466 N8466 N8467 Segment
X8467 N8467 N8468 Segment
X8468 N8468 N8469 Segment
X8469 N8469 N8470 Segment
X8470 N8470 N8471 Segment
X8471 N8471 N8472 Segment
X8472 N8472 N8473 Segment
X8473 N8473 N8474 Segment
X8474 N8474 N8475 Segment
X8475 N8475 N8476 Segment
X8476 N8476 N8477 Segment
X8477 N8477 N8478 Segment
X8478 N8478 N8479 Segment
X8479 N8479 N8480 Segment
X8480 N8480 N8481 Segment
X8481 N8481 N8482 Segment
X8482 N8482 N8483 Segment
X8483 N8483 N8484 Segment
X8484 N8484 N8485 Segment
X8485 N8485 N8486 Segment
X8486 N8486 N8487 Segment
X8487 N8487 N8488 Segment
X8488 N8488 N8489 Segment
X8489 N8489 N8490 Segment
X8490 N8490 N8491 Segment
X8491 N8491 N8492 Segment
X8492 N8492 N8493 Segment
X8493 N8493 N8494 Segment
X8494 N8494 N8495 Segment
X8495 N8495 N8496 Segment
X8496 N8496 N8497 Segment
X8497 N8497 N8498 Segment
X8498 N8498 N8499 Segment
X8499 N8499 N8500 Segment
X8500 N8500 N8501 Segment
X8501 N8501 N8502 Segment
X8502 N8502 N8503 Segment
X8503 N8503 N8504 Segment
X8504 N8504 N8505 Segment
X8505 N8505 N8506 Segment
X8506 N8506 N8507 Segment
X8507 N8507 N8508 Segment
X8508 N8508 N8509 Segment
X8509 N8509 N8510 Segment
X8510 N8510 N8511 Segment
X8511 N8511 N8512 Segment
X8512 N8512 N8513 Segment
X8513 N8513 N8514 Segment
X8514 N8514 N8515 Segment
X8515 N8515 N8516 Segment
X8516 N8516 N8517 Segment
X8517 N8517 N8518 Segment
X8518 N8518 N8519 Segment
X8519 N8519 N8520 Segment
X8520 N8520 N8521 Segment
X8521 N8521 N8522 Segment
X8522 N8522 N8523 Segment
X8523 N8523 N8524 Segment
X8524 N8524 N8525 Segment
X8525 N8525 N8526 Segment
X8526 N8526 N8527 Segment
X8527 N8527 N8528 Segment
X8528 N8528 N8529 Segment
X8529 N8529 N8530 Segment
X8530 N8530 N8531 Segment
X8531 N8531 N8532 Segment
X8532 N8532 N8533 Segment
X8533 N8533 N8534 Segment
X8534 N8534 N8535 Segment
X8535 N8535 N8536 Segment
X8536 N8536 N8537 Segment
X8537 N8537 N8538 Segment
X8538 N8538 N8539 Segment
X8539 N8539 N8540 Segment
X8540 N8540 N8541 Segment
X8541 N8541 N8542 Segment
X8542 N8542 N8543 Segment
X8543 N8543 N8544 Segment
X8544 N8544 N8545 Segment
X8545 N8545 N8546 Segment
X8546 N8546 N8547 Segment
X8547 N8547 N8548 Segment
X8548 N8548 N8549 Segment
X8549 N8549 N8550 Segment
X8550 N8550 N8551 Segment
X8551 N8551 N8552 Segment
X8552 N8552 N8553 Segment
X8553 N8553 N8554 Segment
X8554 N8554 N8555 Segment
X8555 N8555 N8556 Segment
X8556 N8556 N8557 Segment
X8557 N8557 N8558 Segment
X8558 N8558 N8559 Segment
X8559 N8559 N8560 Segment
X8560 N8560 N8561 Segment
X8561 N8561 N8562 Segment
X8562 N8562 N8563 Segment
X8563 N8563 N8564 Segment
X8564 N8564 N8565 Segment
X8565 N8565 N8566 Segment
X8566 N8566 N8567 Segment
X8567 N8567 N8568 Segment
X8568 N8568 N8569 Segment
X8569 N8569 N8570 Segment
X8570 N8570 N8571 Segment
X8571 N8571 N8572 Segment
X8572 N8572 N8573 Segment
X8573 N8573 N8574 Segment
X8574 N8574 N8575 Segment
X8575 N8575 N8576 Segment
X8576 N8576 N8577 Segment
X8577 N8577 N8578 Segment
X8578 N8578 N8579 Segment
X8579 N8579 N8580 Segment
X8580 N8580 N8581 Segment
X8581 N8581 N8582 Segment
X8582 N8582 N8583 Segment
X8583 N8583 N8584 Segment
X8584 N8584 N8585 Segment
X8585 N8585 N8586 Segment
X8586 N8586 N8587 Segment
X8587 N8587 N8588 Segment
X8588 N8588 N8589 Segment
X8589 N8589 N8590 Segment
X8590 N8590 N8591 Segment
X8591 N8591 N8592 Segment
X8592 N8592 N8593 Segment
X8593 N8593 N8594 Segment
X8594 N8594 N8595 Segment
X8595 N8595 N8596 Segment
X8596 N8596 N8597 Segment
X8597 N8597 N8598 Segment
X8598 N8598 N8599 Segment
X8599 N8599 N8600 Segment
X8600 N8600 N8601 Segment
X8601 N8601 N8602 Segment
X8602 N8602 N8603 Segment
X8603 N8603 N8604 Segment
X8604 N8604 N8605 Segment
X8605 N8605 N8606 Segment
X8606 N8606 N8607 Segment
X8607 N8607 N8608 Segment
X8608 N8608 N8609 Segment
X8609 N8609 N8610 Segment
X8610 N8610 N8611 Segment
X8611 N8611 N8612 Segment
X8612 N8612 N8613 Segment
X8613 N8613 N8614 Segment
X8614 N8614 N8615 Segment
X8615 N8615 N8616 Segment
X8616 N8616 N8617 Segment
X8617 N8617 N8618 Segment
X8618 N8618 N8619 Segment
X8619 N8619 N8620 Segment
X8620 N8620 N8621 Segment
X8621 N8621 N8622 Segment
X8622 N8622 N8623 Segment
X8623 N8623 N8624 Segment
X8624 N8624 N8625 Segment
X8625 N8625 N8626 Segment
X8626 N8626 N8627 Segment
X8627 N8627 N8628 Segment
X8628 N8628 N8629 Segment
X8629 N8629 N8630 Segment
X8630 N8630 N8631 Segment
X8631 N8631 N8632 Segment
X8632 N8632 N8633 Segment
X8633 N8633 N8634 Segment
X8634 N8634 N8635 Segment
X8635 N8635 N8636 Segment
X8636 N8636 N8637 Segment
X8637 N8637 N8638 Segment
X8638 N8638 N8639 Segment
X8639 N8639 N8640 Segment
X8640 N8640 N8641 Segment
X8641 N8641 N8642 Segment
X8642 N8642 N8643 Segment
X8643 N8643 N8644 Segment
X8644 N8644 N8645 Segment
X8645 N8645 N8646 Segment
X8646 N8646 N8647 Segment
X8647 N8647 N8648 Segment
X8648 N8648 N8649 Segment
X8649 N8649 N8650 Segment
X8650 N8650 N8651 Segment
X8651 N8651 N8652 Segment
X8652 N8652 N8653 Segment
X8653 N8653 N8654 Segment
X8654 N8654 N8655 Segment
X8655 N8655 N8656 Segment
X8656 N8656 N8657 Segment
X8657 N8657 N8658 Segment
X8658 N8658 N8659 Segment
X8659 N8659 N8660 Segment
X8660 N8660 N8661 Segment
X8661 N8661 N8662 Segment
X8662 N8662 N8663 Segment
X8663 N8663 N8664 Segment
X8664 N8664 N8665 Segment
X8665 N8665 N8666 Segment
X8666 N8666 N8667 Segment
X8667 N8667 N8668 Segment
X8668 N8668 N8669 Segment
X8669 N8669 N8670 Segment
X8670 N8670 N8671 Segment
X8671 N8671 N8672 Segment
X8672 N8672 N8673 Segment
X8673 N8673 N8674 Segment
X8674 N8674 N8675 Segment
X8675 N8675 N8676 Segment
X8676 N8676 N8677 Segment
X8677 N8677 N8678 Segment
X8678 N8678 N8679 Segment
X8679 N8679 N8680 Segment
X8680 N8680 N8681 Segment
X8681 N8681 N8682 Segment
X8682 N8682 N8683 Segment
X8683 N8683 N8684 Segment
X8684 N8684 N8685 Segment
X8685 N8685 N8686 Segment
X8686 N8686 N8687 Segment
X8687 N8687 N8688 Segment
X8688 N8688 N8689 Segment
X8689 N8689 N8690 Segment
X8690 N8690 N8691 Segment
X8691 N8691 N8692 Segment
X8692 N8692 N8693 Segment
X8693 N8693 N8694 Segment
X8694 N8694 N8695 Segment
X8695 N8695 N8696 Segment
X8696 N8696 N8697 Segment
X8697 N8697 N8698 Segment
X8698 N8698 N8699 Segment
X8699 N8699 N8700 Segment
X8700 N8700 N8701 Segment
X8701 N8701 N8702 Segment
X8702 N8702 N8703 Segment
X8703 N8703 N8704 Segment
X8704 N8704 N8705 Segment
X8705 N8705 N8706 Segment
X8706 N8706 N8707 Segment
X8707 N8707 N8708 Segment
X8708 N8708 N8709 Segment
X8709 N8709 N8710 Segment
X8710 N8710 N8711 Segment
X8711 N8711 N8712 Segment
X8712 N8712 N8713 Segment
X8713 N8713 N8714 Segment
X8714 N8714 N8715 Segment
X8715 N8715 N8716 Segment
X8716 N8716 N8717 Segment
X8717 N8717 N8718 Segment
X8718 N8718 N8719 Segment
X8719 N8719 N8720 Segment
X8720 N8720 N8721 Segment
X8721 N8721 N8722 Segment
X8722 N8722 N8723 Segment
X8723 N8723 N8724 Segment
X8724 N8724 N8725 Segment
X8725 N8725 N8726 Segment
X8726 N8726 N8727 Segment
X8727 N8727 N8728 Segment
X8728 N8728 N8729 Segment
X8729 N8729 N8730 Segment
X8730 N8730 N8731 Segment
X8731 N8731 N8732 Segment
X8732 N8732 N8733 Segment
X8733 N8733 N8734 Segment
X8734 N8734 N8735 Segment
X8735 N8735 N8736 Segment
X8736 N8736 N8737 Segment
X8737 N8737 N8738 Segment
X8738 N8738 N8739 Segment
X8739 N8739 N8740 Segment
X8740 N8740 N8741 Segment
X8741 N8741 N8742 Segment
X8742 N8742 N8743 Segment
X8743 N8743 N8744 Segment
X8744 N8744 N8745 Segment
X8745 N8745 N8746 Segment
X8746 N8746 N8747 Segment
X8747 N8747 N8748 Segment
X8748 N8748 N8749 Segment
X8749 N8749 N8750 Segment
X8750 N8750 N8751 Segment
X8751 N8751 N8752 Segment
X8752 N8752 N8753 Segment
X8753 N8753 N8754 Segment
X8754 N8754 N8755 Segment
X8755 N8755 N8756 Segment
X8756 N8756 N8757 Segment
X8757 N8757 N8758 Segment
X8758 N8758 N8759 Segment
X8759 N8759 N8760 Segment
X8760 N8760 N8761 Segment
X8761 N8761 N8762 Segment
X8762 N8762 N8763 Segment
X8763 N8763 N8764 Segment
X8764 N8764 N8765 Segment
X8765 N8765 N8766 Segment
X8766 N8766 N8767 Segment
X8767 N8767 N8768 Segment
X8768 N8768 N8769 Segment
X8769 N8769 N8770 Segment
X8770 N8770 N8771 Segment
X8771 N8771 N8772 Segment
X8772 N8772 N8773 Segment
X8773 N8773 N8774 Segment
X8774 N8774 N8775 Segment
X8775 N8775 N8776 Segment
X8776 N8776 N8777 Segment
X8777 N8777 N8778 Segment
X8778 N8778 N8779 Segment
X8779 N8779 N8780 Segment
X8780 N8780 N8781 Segment
X8781 N8781 N8782 Segment
X8782 N8782 N8783 Segment
X8783 N8783 N8784 Segment
X8784 N8784 N8785 Segment
X8785 N8785 N8786 Segment
X8786 N8786 N8787 Segment
X8787 N8787 N8788 Segment
X8788 N8788 N8789 Segment
X8789 N8789 N8790 Segment
X8790 N8790 N8791 Segment
X8791 N8791 N8792 Segment
X8792 N8792 N8793 Segment
X8793 N8793 N8794 Segment
X8794 N8794 N8795 Segment
X8795 N8795 N8796 Segment
X8796 N8796 N8797 Segment
X8797 N8797 N8798 Segment
X8798 N8798 N8799 Segment
X8799 N8799 N8800 Segment
X8800 N8800 N8801 Segment
X8801 N8801 N8802 Segment
X8802 N8802 N8803 Segment
X8803 N8803 N8804 Segment
X8804 N8804 N8805 Segment
X8805 N8805 N8806 Segment
X8806 N8806 N8807 Segment
X8807 N8807 N8808 Segment
X8808 N8808 N8809 Segment
X8809 N8809 N8810 Segment
X8810 N8810 N8811 Segment
X8811 N8811 N8812 Segment
X8812 N8812 N8813 Segment
X8813 N8813 N8814 Segment
X8814 N8814 N8815 Segment
X8815 N8815 N8816 Segment
X8816 N8816 N8817 Segment
X8817 N8817 N8818 Segment
X8818 N8818 N8819 Segment
X8819 N8819 N8820 Segment
X8820 N8820 N8821 Segment
X8821 N8821 N8822 Segment
X8822 N8822 N8823 Segment
X8823 N8823 N8824 Segment
X8824 N8824 N8825 Segment
X8825 N8825 N8826 Segment
X8826 N8826 N8827 Segment
X8827 N8827 N8828 Segment
X8828 N8828 N8829 Segment
X8829 N8829 N8830 Segment
X8830 N8830 N8831 Segment
X8831 N8831 N8832 Segment
X8832 N8832 N8833 Segment
X8833 N8833 N8834 Segment
X8834 N8834 N8835 Segment
X8835 N8835 N8836 Segment
X8836 N8836 N8837 Segment
X8837 N8837 N8838 Segment
X8838 N8838 N8839 Segment
X8839 N8839 N8840 Segment
X8840 N8840 N8841 Segment
X8841 N8841 N8842 Segment
X8842 N8842 N8843 Segment
X8843 N8843 N8844 Segment
X8844 N8844 N8845 Segment
X8845 N8845 N8846 Segment
X8846 N8846 N8847 Segment
X8847 N8847 N8848 Segment
X8848 N8848 N8849 Segment
X8849 N8849 N8850 Segment
X8850 N8850 N8851 Segment
X8851 N8851 N8852 Segment
X8852 N8852 N8853 Segment
X8853 N8853 N8854 Segment
X8854 N8854 N8855 Segment
X8855 N8855 N8856 Segment
X8856 N8856 N8857 Segment
X8857 N8857 N8858 Segment
X8858 N8858 N8859 Segment
X8859 N8859 N8860 Segment
X8860 N8860 N8861 Segment
X8861 N8861 N8862 Segment
X8862 N8862 N8863 Segment
X8863 N8863 N8864 Segment
X8864 N8864 N8865 Segment
X8865 N8865 N8866 Segment
X8866 N8866 N8867 Segment
X8867 N8867 N8868 Segment
X8868 N8868 N8869 Segment
X8869 N8869 N8870 Segment
X8870 N8870 N8871 Segment
X8871 N8871 N8872 Segment
X8872 N8872 N8873 Segment
X8873 N8873 N8874 Segment
X8874 N8874 N8875 Segment
X8875 N8875 N8876 Segment
X8876 N8876 N8877 Segment
X8877 N8877 N8878 Segment
X8878 N8878 N8879 Segment
X8879 N8879 N8880 Segment
X8880 N8880 N8881 Segment
X8881 N8881 N8882 Segment
X8882 N8882 N8883 Segment
X8883 N8883 N8884 Segment
X8884 N8884 N8885 Segment
X8885 N8885 N8886 Segment
X8886 N8886 N8887 Segment
X8887 N8887 N8888 Segment
X8888 N8888 N8889 Segment
X8889 N8889 N8890 Segment
X8890 N8890 N8891 Segment
X8891 N8891 N8892 Segment
X8892 N8892 N8893 Segment
X8893 N8893 N8894 Segment
X8894 N8894 N8895 Segment
X8895 N8895 N8896 Segment
X8896 N8896 N8897 Segment
X8897 N8897 N8898 Segment
X8898 N8898 N8899 Segment
X8899 N8899 N8900 Segment
X8900 N8900 N8901 Segment
X8901 N8901 N8902 Segment
X8902 N8902 N8903 Segment
X8903 N8903 N8904 Segment
X8904 N8904 N8905 Segment
X8905 N8905 N8906 Segment
X8906 N8906 N8907 Segment
X8907 N8907 N8908 Segment
X8908 N8908 N8909 Segment
X8909 N8909 N8910 Segment
X8910 N8910 N8911 Segment
X8911 N8911 N8912 Segment
X8912 N8912 N8913 Segment
X8913 N8913 N8914 Segment
X8914 N8914 N8915 Segment
X8915 N8915 N8916 Segment
X8916 N8916 N8917 Segment
X8917 N8917 N8918 Segment
X8918 N8918 N8919 Segment
X8919 N8919 N8920 Segment
X8920 N8920 N8921 Segment
X8921 N8921 N8922 Segment
X8922 N8922 N8923 Segment
X8923 N8923 N8924 Segment
X8924 N8924 N8925 Segment
X8925 N8925 N8926 Segment
X8926 N8926 N8927 Segment
X8927 N8927 N8928 Segment
X8928 N8928 N8929 Segment
X8929 N8929 N8930 Segment
X8930 N8930 N8931 Segment
X8931 N8931 N8932 Segment
X8932 N8932 N8933 Segment
X8933 N8933 N8934 Segment
X8934 N8934 N8935 Segment
X8935 N8935 N8936 Segment
X8936 N8936 N8937 Segment
X8937 N8937 N8938 Segment
X8938 N8938 N8939 Segment
X8939 N8939 N8940 Segment
X8940 N8940 N8941 Segment
X8941 N8941 N8942 Segment
X8942 N8942 N8943 Segment
X8943 N8943 N8944 Segment
X8944 N8944 N8945 Segment
X8945 N8945 N8946 Segment
X8946 N8946 N8947 Segment
X8947 N8947 N8948 Segment
X8948 N8948 N8949 Segment
X8949 N8949 N8950 Segment
X8950 N8950 N8951 Segment
X8951 N8951 N8952 Segment
X8952 N8952 N8953 Segment
X8953 N8953 N8954 Segment
X8954 N8954 N8955 Segment
X8955 N8955 N8956 Segment
X8956 N8956 N8957 Segment
X8957 N8957 N8958 Segment
X8958 N8958 N8959 Segment
X8959 N8959 N8960 Segment
X8960 N8960 N8961 Segment
X8961 N8961 N8962 Segment
X8962 N8962 N8963 Segment
X8963 N8963 N8964 Segment
X8964 N8964 N8965 Segment
X8965 N8965 N8966 Segment
X8966 N8966 N8967 Segment
X8967 N8967 N8968 Segment
X8968 N8968 N8969 Segment
X8969 N8969 N8970 Segment
X8970 N8970 N8971 Segment
X8971 N8971 N8972 Segment
X8972 N8972 N8973 Segment
X8973 N8973 N8974 Segment
X8974 N8974 N8975 Segment
X8975 N8975 N8976 Segment
X8976 N8976 N8977 Segment
X8977 N8977 N8978 Segment
X8978 N8978 N8979 Segment
X8979 N8979 N8980 Segment
X8980 N8980 N8981 Segment
X8981 N8981 N8982 Segment
X8982 N8982 N8983 Segment
X8983 N8983 N8984 Segment
X8984 N8984 N8985 Segment
X8985 N8985 N8986 Segment
X8986 N8986 N8987 Segment
X8987 N8987 N8988 Segment
X8988 N8988 N8989 Segment
X8989 N8989 N8990 Segment
X8990 N8990 N8991 Segment
X8991 N8991 N8992 Segment
X8992 N8992 N8993 Segment
X8993 N8993 N8994 Segment
X8994 N8994 N8995 Segment
X8995 N8995 N8996 Segment
X8996 N8996 N8997 Segment
X8997 N8997 N8998 Segment
X8998 N8998 N8999 Segment
X8999 N8999 N9000 Segment
X9000 N9000 N9001 Segment
X9001 N9001 N9002 Segment
X9002 N9002 N9003 Segment
X9003 N9003 N9004 Segment
X9004 N9004 N9005 Segment
X9005 N9005 N9006 Segment
X9006 N9006 N9007 Segment
X9007 N9007 N9008 Segment
X9008 N9008 N9009 Segment
X9009 N9009 N9010 Segment
X9010 N9010 N9011 Segment
X9011 N9011 N9012 Segment
X9012 N9012 N9013 Segment
X9013 N9013 N9014 Segment
X9014 N9014 N9015 Segment
X9015 N9015 N9016 Segment
X9016 N9016 N9017 Segment
X9017 N9017 N9018 Segment
X9018 N9018 N9019 Segment
X9019 N9019 N9020 Segment
X9020 N9020 N9021 Segment
X9021 N9021 N9022 Segment
X9022 N9022 N9023 Segment
X9023 N9023 N9024 Segment
X9024 N9024 N9025 Segment
X9025 N9025 N9026 Segment
X9026 N9026 N9027 Segment
X9027 N9027 N9028 Segment
X9028 N9028 N9029 Segment
X9029 N9029 N9030 Segment
X9030 N9030 N9031 Segment
X9031 N9031 N9032 Segment
X9032 N9032 N9033 Segment
X9033 N9033 N9034 Segment
X9034 N9034 N9035 Segment
X9035 N9035 N9036 Segment
X9036 N9036 N9037 Segment
X9037 N9037 N9038 Segment
X9038 N9038 N9039 Segment
X9039 N9039 N9040 Segment
X9040 N9040 N9041 Segment
X9041 N9041 N9042 Segment
X9042 N9042 N9043 Segment
X9043 N9043 N9044 Segment
X9044 N9044 N9045 Segment
X9045 N9045 N9046 Segment
X9046 N9046 N9047 Segment
X9047 N9047 N9048 Segment
X9048 N9048 N9049 Segment
X9049 N9049 N9050 Segment
X9050 N9050 N9051 Segment
X9051 N9051 N9052 Segment
X9052 N9052 N9053 Segment
X9053 N9053 N9054 Segment
X9054 N9054 N9055 Segment
X9055 N9055 N9056 Segment
X9056 N9056 N9057 Segment
X9057 N9057 N9058 Segment
X9058 N9058 N9059 Segment
X9059 N9059 N9060 Segment
X9060 N9060 N9061 Segment
X9061 N9061 N9062 Segment
X9062 N9062 N9063 Segment
X9063 N9063 N9064 Segment
X9064 N9064 N9065 Segment
X9065 N9065 N9066 Segment
X9066 N9066 N9067 Segment
X9067 N9067 N9068 Segment
X9068 N9068 N9069 Segment
X9069 N9069 N9070 Segment
X9070 N9070 N9071 Segment
X9071 N9071 N9072 Segment
X9072 N9072 N9073 Segment
X9073 N9073 N9074 Segment
X9074 N9074 N9075 Segment
X9075 N9075 N9076 Segment
X9076 N9076 N9077 Segment
X9077 N9077 N9078 Segment
X9078 N9078 N9079 Segment
X9079 N9079 N9080 Segment
X9080 N9080 N9081 Segment
X9081 N9081 N9082 Segment
X9082 N9082 N9083 Segment
X9083 N9083 N9084 Segment
X9084 N9084 N9085 Segment
X9085 N9085 N9086 Segment
X9086 N9086 N9087 Segment
X9087 N9087 N9088 Segment
X9088 N9088 N9089 Segment
X9089 N9089 N9090 Segment
X9090 N9090 N9091 Segment
X9091 N9091 N9092 Segment
X9092 N9092 N9093 Segment
X9093 N9093 N9094 Segment
X9094 N9094 N9095 Segment
X9095 N9095 N9096 Segment
X9096 N9096 N9097 Segment
X9097 N9097 N9098 Segment
X9098 N9098 N9099 Segment
X9099 N9099 N9100 Segment
X9100 N9100 N9101 Segment
X9101 N9101 N9102 Segment
X9102 N9102 N9103 Segment
X9103 N9103 N9104 Segment
X9104 N9104 N9105 Segment
X9105 N9105 N9106 Segment
X9106 N9106 N9107 Segment
X9107 N9107 N9108 Segment
X9108 N9108 N9109 Segment
X9109 N9109 N9110 Segment
X9110 N9110 N9111 Segment
X9111 N9111 N9112 Segment
X9112 N9112 N9113 Segment
X9113 N9113 N9114 Segment
X9114 N9114 N9115 Segment
X9115 N9115 N9116 Segment
X9116 N9116 N9117 Segment
X9117 N9117 N9118 Segment
X9118 N9118 N9119 Segment
X9119 N9119 N9120 Segment
X9120 N9120 N9121 Segment
X9121 N9121 N9122 Segment
X9122 N9122 N9123 Segment
X9123 N9123 N9124 Segment
X9124 N9124 N9125 Segment
X9125 N9125 N9126 Segment
X9126 N9126 N9127 Segment
X9127 N9127 N9128 Segment
X9128 N9128 N9129 Segment
X9129 N9129 N9130 Segment
X9130 N9130 N9131 Segment
X9131 N9131 N9132 Segment
X9132 N9132 N9133 Segment
X9133 N9133 N9134 Segment
X9134 N9134 N9135 Segment
X9135 N9135 N9136 Segment
X9136 N9136 N9137 Segment
X9137 N9137 N9138 Segment
X9138 N9138 N9139 Segment
X9139 N9139 N9140 Segment
X9140 N9140 N9141 Segment
X9141 N9141 N9142 Segment
X9142 N9142 N9143 Segment
X9143 N9143 N9144 Segment
X9144 N9144 N9145 Segment
X9145 N9145 N9146 Segment
X9146 N9146 N9147 Segment
X9147 N9147 N9148 Segment
X9148 N9148 N9149 Segment
X9149 N9149 N9150 Segment
X9150 N9150 N9151 Segment
X9151 N9151 N9152 Segment
X9152 N9152 N9153 Segment
X9153 N9153 N9154 Segment
X9154 N9154 N9155 Segment
X9155 N9155 N9156 Segment
X9156 N9156 N9157 Segment
X9157 N9157 N9158 Segment
X9158 N9158 N9159 Segment
X9159 N9159 N9160 Segment
X9160 N9160 N9161 Segment
X9161 N9161 N9162 Segment
X9162 N9162 N9163 Segment
X9163 N9163 N9164 Segment
X9164 N9164 N9165 Segment
X9165 N9165 N9166 Segment
X9166 N9166 N9167 Segment
X9167 N9167 N9168 Segment
X9168 N9168 N9169 Segment
X9169 N9169 N9170 Segment
X9170 N9170 N9171 Segment
X9171 N9171 N9172 Segment
X9172 N9172 N9173 Segment
X9173 N9173 N9174 Segment
X9174 N9174 N9175 Segment
X9175 N9175 N9176 Segment
X9176 N9176 N9177 Segment
X9177 N9177 N9178 Segment
X9178 N9178 N9179 Segment
X9179 N9179 N9180 Segment
X9180 N9180 N9181 Segment
X9181 N9181 N9182 Segment
X9182 N9182 N9183 Segment
X9183 N9183 N9184 Segment
X9184 N9184 N9185 Segment
X9185 N9185 N9186 Segment
X9186 N9186 N9187 Segment
X9187 N9187 N9188 Segment
X9188 N9188 N9189 Segment
X9189 N9189 N9190 Segment
X9190 N9190 N9191 Segment
X9191 N9191 N9192 Segment
X9192 N9192 N9193 Segment
X9193 N9193 N9194 Segment
X9194 N9194 N9195 Segment
X9195 N9195 N9196 Segment
X9196 N9196 N9197 Segment
X9197 N9197 N9198 Segment
X9198 N9198 N9199 Segment
X9199 N9199 N9200 Segment
X9200 N9200 N9201 Segment
X9201 N9201 N9202 Segment
X9202 N9202 N9203 Segment
X9203 N9203 N9204 Segment
X9204 N9204 N9205 Segment
X9205 N9205 N9206 Segment
X9206 N9206 N9207 Segment
X9207 N9207 N9208 Segment
X9208 N9208 N9209 Segment
X9209 N9209 N9210 Segment
X9210 N9210 N9211 Segment
X9211 N9211 N9212 Segment
X9212 N9212 N9213 Segment
X9213 N9213 N9214 Segment
X9214 N9214 N9215 Segment
X9215 N9215 N9216 Segment
X9216 N9216 N9217 Segment
X9217 N9217 N9218 Segment
X9218 N9218 N9219 Segment
X9219 N9219 N9220 Segment
X9220 N9220 N9221 Segment
X9221 N9221 N9222 Segment
X9222 N9222 N9223 Segment
X9223 N9223 N9224 Segment
X9224 N9224 N9225 Segment
X9225 N9225 N9226 Segment
X9226 N9226 N9227 Segment
X9227 N9227 N9228 Segment
X9228 N9228 N9229 Segment
X9229 N9229 N9230 Segment
X9230 N9230 N9231 Segment
X9231 N9231 N9232 Segment
X9232 N9232 N9233 Segment
X9233 N9233 N9234 Segment
X9234 N9234 N9235 Segment
X9235 N9235 N9236 Segment
X9236 N9236 N9237 Segment
X9237 N9237 N9238 Segment
X9238 N9238 N9239 Segment
X9239 N9239 N9240 Segment
X9240 N9240 N9241 Segment
X9241 N9241 N9242 Segment
X9242 N9242 N9243 Segment
X9243 N9243 N9244 Segment
X9244 N9244 N9245 Segment
X9245 N9245 N9246 Segment
X9246 N9246 N9247 Segment
X9247 N9247 N9248 Segment
X9248 N9248 N9249 Segment
X9249 N9249 N9250 Segment
X9250 N9250 N9251 Segment
X9251 N9251 N9252 Segment
X9252 N9252 N9253 Segment
X9253 N9253 N9254 Segment
X9254 N9254 N9255 Segment
X9255 N9255 N9256 Segment
X9256 N9256 N9257 Segment
X9257 N9257 N9258 Segment
X9258 N9258 N9259 Segment
X9259 N9259 N9260 Segment
X9260 N9260 N9261 Segment
X9261 N9261 N9262 Segment
X9262 N9262 N9263 Segment
X9263 N9263 N9264 Segment
X9264 N9264 N9265 Segment
X9265 N9265 N9266 Segment
X9266 N9266 N9267 Segment
X9267 N9267 N9268 Segment
X9268 N9268 N9269 Segment
X9269 N9269 N9270 Segment
X9270 N9270 N9271 Segment
X9271 N9271 N9272 Segment
X9272 N9272 N9273 Segment
X9273 N9273 N9274 Segment
X9274 N9274 N9275 Segment
X9275 N9275 N9276 Segment
X9276 N9276 N9277 Segment
X9277 N9277 N9278 Segment
X9278 N9278 N9279 Segment
X9279 N9279 N9280 Segment
X9280 N9280 N9281 Segment
X9281 N9281 N9282 Segment
X9282 N9282 N9283 Segment
X9283 N9283 N9284 Segment
X9284 N9284 N9285 Segment
X9285 N9285 N9286 Segment
X9286 N9286 N9287 Segment
X9287 N9287 N9288 Segment
X9288 N9288 N9289 Segment
X9289 N9289 N9290 Segment
X9290 N9290 N9291 Segment
X9291 N9291 N9292 Segment
X9292 N9292 N9293 Segment
X9293 N9293 N9294 Segment
X9294 N9294 N9295 Segment
X9295 N9295 N9296 Segment
X9296 N9296 N9297 Segment
X9297 N9297 N9298 Segment
X9298 N9298 N9299 Segment
X9299 N9299 N9300 Segment
X9300 N9300 N9301 Segment
X9301 N9301 N9302 Segment
X9302 N9302 N9303 Segment
X9303 N9303 N9304 Segment
X9304 N9304 N9305 Segment
X9305 N9305 N9306 Segment
X9306 N9306 N9307 Segment
X9307 N9307 N9308 Segment
X9308 N9308 N9309 Segment
X9309 N9309 N9310 Segment
X9310 N9310 N9311 Segment
X9311 N9311 N9312 Segment
X9312 N9312 N9313 Segment
X9313 N9313 N9314 Segment
X9314 N9314 N9315 Segment
X9315 N9315 N9316 Segment
X9316 N9316 N9317 Segment
X9317 N9317 N9318 Segment
X9318 N9318 N9319 Segment
X9319 N9319 N9320 Segment
X9320 N9320 N9321 Segment
X9321 N9321 N9322 Segment
X9322 N9322 N9323 Segment
X9323 N9323 N9324 Segment
X9324 N9324 N9325 Segment
X9325 N9325 N9326 Segment
X9326 N9326 N9327 Segment
X9327 N9327 N9328 Segment
X9328 N9328 N9329 Segment
X9329 N9329 N9330 Segment
X9330 N9330 N9331 Segment
X9331 N9331 N9332 Segment
X9332 N9332 N9333 Segment
X9333 N9333 N9334 Segment
X9334 N9334 N9335 Segment
X9335 N9335 N9336 Segment
X9336 N9336 N9337 Segment
X9337 N9337 N9338 Segment
X9338 N9338 N9339 Segment
X9339 N9339 N9340 Segment
X9340 N9340 N9341 Segment
X9341 N9341 N9342 Segment
X9342 N9342 N9343 Segment
X9343 N9343 N9344 Segment
X9344 N9344 N9345 Segment
X9345 N9345 N9346 Segment
X9346 N9346 N9347 Segment
X9347 N9347 N9348 Segment
X9348 N9348 N9349 Segment
X9349 N9349 N9350 Segment
X9350 N9350 N9351 Segment
X9351 N9351 N9352 Segment
X9352 N9352 N9353 Segment
X9353 N9353 N9354 Segment
X9354 N9354 N9355 Segment
X9355 N9355 N9356 Segment
X9356 N9356 N9357 Segment
X9357 N9357 N9358 Segment
X9358 N9358 N9359 Segment
X9359 N9359 N9360 Segment
X9360 N9360 N9361 Segment
X9361 N9361 N9362 Segment
X9362 N9362 N9363 Segment
X9363 N9363 N9364 Segment
X9364 N9364 N9365 Segment
X9365 N9365 N9366 Segment
X9366 N9366 N9367 Segment
X9367 N9367 N9368 Segment
X9368 N9368 N9369 Segment
X9369 N9369 N9370 Segment
X9370 N9370 N9371 Segment
X9371 N9371 N9372 Segment
X9372 N9372 N9373 Segment
X9373 N9373 N9374 Segment
X9374 N9374 N9375 Segment
X9375 N9375 N9376 Segment
X9376 N9376 N9377 Segment
X9377 N9377 N9378 Segment
X9378 N9378 N9379 Segment
X9379 N9379 N9380 Segment
X9380 N9380 N9381 Segment
X9381 N9381 N9382 Segment
X9382 N9382 N9383 Segment
X9383 N9383 N9384 Segment
X9384 N9384 N9385 Segment
X9385 N9385 N9386 Segment
X9386 N9386 N9387 Segment
X9387 N9387 N9388 Segment
X9388 N9388 N9389 Segment
X9389 N9389 N9390 Segment
X9390 N9390 N9391 Segment
X9391 N9391 N9392 Segment
X9392 N9392 N9393 Segment
X9393 N9393 N9394 Segment
X9394 N9394 N9395 Segment
X9395 N9395 N9396 Segment
X9396 N9396 N9397 Segment
X9397 N9397 N9398 Segment
X9398 N9398 N9399 Segment
X9399 N9399 N9400 Segment
X9400 N9400 N9401 Segment
X9401 N9401 N9402 Segment
X9402 N9402 N9403 Segment
X9403 N9403 N9404 Segment
X9404 N9404 N9405 Segment
X9405 N9405 N9406 Segment
X9406 N9406 N9407 Segment
X9407 N9407 N9408 Segment
X9408 N9408 N9409 Segment
X9409 N9409 N9410 Segment
X9410 N9410 N9411 Segment
X9411 N9411 N9412 Segment
X9412 N9412 N9413 Segment
X9413 N9413 N9414 Segment
X9414 N9414 N9415 Segment
X9415 N9415 N9416 Segment
X9416 N9416 N9417 Segment
X9417 N9417 N9418 Segment
X9418 N9418 N9419 Segment
X9419 N9419 N9420 Segment
X9420 N9420 N9421 Segment
X9421 N9421 N9422 Segment
X9422 N9422 N9423 Segment
X9423 N9423 N9424 Segment
X9424 N9424 N9425 Segment
X9425 N9425 N9426 Segment
X9426 N9426 N9427 Segment
X9427 N9427 N9428 Segment
X9428 N9428 N9429 Segment
X9429 N9429 N9430 Segment
X9430 N9430 N9431 Segment
X9431 N9431 N9432 Segment
X9432 N9432 N9433 Segment
X9433 N9433 N9434 Segment
X9434 N9434 N9435 Segment
X9435 N9435 N9436 Segment
X9436 N9436 N9437 Segment
X9437 N9437 N9438 Segment
X9438 N9438 N9439 Segment
X9439 N9439 N9440 Segment
X9440 N9440 N9441 Segment
X9441 N9441 N9442 Segment
X9442 N9442 N9443 Segment
X9443 N9443 N9444 Segment
X9444 N9444 N9445 Segment
X9445 N9445 N9446 Segment
X9446 N9446 N9447 Segment
X9447 N9447 N9448 Segment
X9448 N9448 N9449 Segment
X9449 N9449 N9450 Segment
X9450 N9450 N9451 Segment
X9451 N9451 N9452 Segment
X9452 N9452 N9453 Segment
X9453 N9453 N9454 Segment
X9454 N9454 N9455 Segment
X9455 N9455 N9456 Segment
X9456 N9456 N9457 Segment
X9457 N9457 N9458 Segment
X9458 N9458 N9459 Segment
X9459 N9459 N9460 Segment
X9460 N9460 N9461 Segment
X9461 N9461 N9462 Segment
X9462 N9462 N9463 Segment
X9463 N9463 N9464 Segment
X9464 N9464 N9465 Segment
X9465 N9465 N9466 Segment
X9466 N9466 N9467 Segment
X9467 N9467 N9468 Segment
X9468 N9468 N9469 Segment
X9469 N9469 N9470 Segment
X9470 N9470 N9471 Segment
X9471 N9471 N9472 Segment
X9472 N9472 N9473 Segment
X9473 N9473 N9474 Segment
X9474 N9474 N9475 Segment
X9475 N9475 N9476 Segment
X9476 N9476 N9477 Segment
X9477 N9477 N9478 Segment
X9478 N9478 N9479 Segment
X9479 N9479 N9480 Segment
X9480 N9480 N9481 Segment
X9481 N9481 N9482 Segment
X9482 N9482 N9483 Segment
X9483 N9483 N9484 Segment
X9484 N9484 N9485 Segment
X9485 N9485 N9486 Segment
X9486 N9486 N9487 Segment
X9487 N9487 N9488 Segment
X9488 N9488 N9489 Segment
X9489 N9489 N9490 Segment
X9490 N9490 N9491 Segment
X9491 N9491 N9492 Segment
X9492 N9492 N9493 Segment
X9493 N9493 N9494 Segment
X9494 N9494 N9495 Segment
X9495 N9495 N9496 Segment
X9496 N9496 N9497 Segment
X9497 N9497 N9498 Segment
X9498 N9498 N9499 Segment
X9499 N9499 N9500 Segment
X9500 N9500 N9501 Segment
X9501 N9501 N9502 Segment
X9502 N9502 N9503 Segment
X9503 N9503 N9504 Segment
X9504 N9504 N9505 Segment
X9505 N9505 N9506 Segment
X9506 N9506 N9507 Segment
X9507 N9507 N9508 Segment
X9508 N9508 N9509 Segment
X9509 N9509 N9510 Segment
X9510 N9510 N9511 Segment
X9511 N9511 N9512 Segment
X9512 N9512 N9513 Segment
X9513 N9513 N9514 Segment
X9514 N9514 N9515 Segment
X9515 N9515 N9516 Segment
X9516 N9516 N9517 Segment
X9517 N9517 N9518 Segment
X9518 N9518 N9519 Segment
X9519 N9519 N9520 Segment
X9520 N9520 N9521 Segment
X9521 N9521 N9522 Segment
X9522 N9522 N9523 Segment
X9523 N9523 N9524 Segment
X9524 N9524 N9525 Segment
X9525 N9525 N9526 Segment
X9526 N9526 N9527 Segment
X9527 N9527 N9528 Segment
X9528 N9528 N9529 Segment
X9529 N9529 N9530 Segment
X9530 N9530 N9531 Segment
X9531 N9531 N9532 Segment
X9532 N9532 N9533 Segment
X9533 N9533 N9534 Segment
X9534 N9534 N9535 Segment
X9535 N9535 N9536 Segment
X9536 N9536 N9537 Segment
X9537 N9537 N9538 Segment
X9538 N9538 N9539 Segment
X9539 N9539 N9540 Segment
X9540 N9540 N9541 Segment
X9541 N9541 N9542 Segment
X9542 N9542 N9543 Segment
X9543 N9543 N9544 Segment
X9544 N9544 N9545 Segment
X9545 N9545 N9546 Segment
X9546 N9546 N9547 Segment
X9547 N9547 N9548 Segment
X9548 N9548 N9549 Segment
X9549 N9549 N9550 Segment
X9550 N9550 N9551 Segment
X9551 N9551 N9552 Segment
X9552 N9552 N9553 Segment
X9553 N9553 N9554 Segment
X9554 N9554 N9555 Segment
X9555 N9555 N9556 Segment
X9556 N9556 N9557 Segment
X9557 N9557 N9558 Segment
X9558 N9558 N9559 Segment
X9559 N9559 N9560 Segment
X9560 N9560 N9561 Segment
X9561 N9561 N9562 Segment
X9562 N9562 N9563 Segment
X9563 N9563 N9564 Segment
X9564 N9564 N9565 Segment
X9565 N9565 N9566 Segment
X9566 N9566 N9567 Segment
X9567 N9567 N9568 Segment
X9568 N9568 N9569 Segment
X9569 N9569 N9570 Segment
X9570 N9570 N9571 Segment
X9571 N9571 N9572 Segment
X9572 N9572 N9573 Segment
X9573 N9573 N9574 Segment
X9574 N9574 N9575 Segment
X9575 N9575 N9576 Segment
X9576 N9576 N9577 Segment
X9577 N9577 N9578 Segment
X9578 N9578 N9579 Segment
X9579 N9579 N9580 Segment
X9580 N9580 N9581 Segment
X9581 N9581 N9582 Segment
X9582 N9582 N9583 Segment
X9583 N9583 N9584 Segment
X9584 N9584 N9585 Segment
X9585 N9585 N9586 Segment
X9586 N9586 N9587 Segment
X9587 N9587 N9588 Segment
X9588 N9588 N9589 Segment
X9589 N9589 N9590 Segment
X9590 N9590 N9591 Segment
X9591 N9591 N9592 Segment
X9592 N9592 N9593 Segment
X9593 N9593 N9594 Segment
X9594 N9594 N9595 Segment
X9595 N9595 N9596 Segment
X9596 N9596 N9597 Segment
X9597 N9597 N9598 Segment
X9598 N9598 N9599 Segment
X9599 N9599 N9600 Segment
X9600 N9600 N9601 Segment
X9601 N9601 N9602 Segment
X9602 N9602 N9603 Segment
X9603 N9603 N9604 Segment
X9604 N9604 N9605 Segment
X9605 N9605 N9606 Segment
X9606 N9606 N9607 Segment
X9607 N9607 N9608 Segment
X9608 N9608 N9609 Segment
X9609 N9609 N9610 Segment
X9610 N9610 N9611 Segment
X9611 N9611 N9612 Segment
X9612 N9612 N9613 Segment
X9613 N9613 N9614 Segment
X9614 N9614 N9615 Segment
X9615 N9615 N9616 Segment
X9616 N9616 N9617 Segment
X9617 N9617 N9618 Segment
X9618 N9618 N9619 Segment
X9619 N9619 N9620 Segment
X9620 N9620 N9621 Segment
X9621 N9621 N9622 Segment
X9622 N9622 N9623 Segment
X9623 N9623 N9624 Segment
X9624 N9624 N9625 Segment
X9625 N9625 N9626 Segment
X9626 N9626 N9627 Segment
X9627 N9627 N9628 Segment
X9628 N9628 N9629 Segment
X9629 N9629 N9630 Segment
X9630 N9630 N9631 Segment
X9631 N9631 N9632 Segment
X9632 N9632 N9633 Segment
X9633 N9633 N9634 Segment
X9634 N9634 N9635 Segment
X9635 N9635 N9636 Segment
X9636 N9636 N9637 Segment
X9637 N9637 N9638 Segment
X9638 N9638 N9639 Segment
X9639 N9639 N9640 Segment
X9640 N9640 N9641 Segment
X9641 N9641 N9642 Segment
X9642 N9642 N9643 Segment
X9643 N9643 N9644 Segment
X9644 N9644 N9645 Segment
X9645 N9645 N9646 Segment
X9646 N9646 N9647 Segment
X9647 N9647 N9648 Segment
X9648 N9648 N9649 Segment
X9649 N9649 N9650 Segment
X9650 N9650 N9651 Segment
X9651 N9651 N9652 Segment
X9652 N9652 N9653 Segment
X9653 N9653 N9654 Segment
X9654 N9654 N9655 Segment
X9655 N9655 N9656 Segment
X9656 N9656 N9657 Segment
X9657 N9657 N9658 Segment
X9658 N9658 N9659 Segment
X9659 N9659 N9660 Segment
X9660 N9660 N9661 Segment
X9661 N9661 N9662 Segment
X9662 N9662 N9663 Segment
X9663 N9663 N9664 Segment
X9664 N9664 N9665 Segment
X9665 N9665 N9666 Segment
X9666 N9666 N9667 Segment
X9667 N9667 N9668 Segment
X9668 N9668 N9669 Segment
X9669 N9669 N9670 Segment
X9670 N9670 N9671 Segment
X9671 N9671 N9672 Segment
X9672 N9672 N9673 Segment
X9673 N9673 N9674 Segment
X9674 N9674 N9675 Segment
X9675 N9675 N9676 Segment
X9676 N9676 N9677 Segment
X9677 N9677 N9678 Segment
X9678 N9678 N9679 Segment
X9679 N9679 N9680 Segment
X9680 N9680 N9681 Segment
X9681 N9681 N9682 Segment
X9682 N9682 N9683 Segment
X9683 N9683 N9684 Segment
X9684 N9684 N9685 Segment
X9685 N9685 N9686 Segment
X9686 N9686 N9687 Segment
X9687 N9687 N9688 Segment
X9688 N9688 N9689 Segment
X9689 N9689 N9690 Segment
X9690 N9690 N9691 Segment
X9691 N9691 N9692 Segment
X9692 N9692 N9693 Segment
X9693 N9693 N9694 Segment
X9694 N9694 N9695 Segment
X9695 N9695 N9696 Segment
X9696 N9696 N9697 Segment
X9697 N9697 N9698 Segment
X9698 N9698 N9699 Segment
X9699 N9699 N9700 Segment
X9700 N9700 N9701 Segment
X9701 N9701 N9702 Segment
X9702 N9702 N9703 Segment
X9703 N9703 N9704 Segment
X9704 N9704 N9705 Segment
X9705 N9705 N9706 Segment
X9706 N9706 N9707 Segment
X9707 N9707 N9708 Segment
X9708 N9708 N9709 Segment
X9709 N9709 N9710 Segment
X9710 N9710 N9711 Segment
X9711 N9711 N9712 Segment
X9712 N9712 N9713 Segment
X9713 N9713 N9714 Segment
X9714 N9714 N9715 Segment
X9715 N9715 N9716 Segment
X9716 N9716 N9717 Segment
X9717 N9717 N9718 Segment
X9718 N9718 N9719 Segment
X9719 N9719 N9720 Segment
X9720 N9720 N9721 Segment
X9721 N9721 N9722 Segment
X9722 N9722 N9723 Segment
X9723 N9723 N9724 Segment
X9724 N9724 N9725 Segment
X9725 N9725 N9726 Segment
X9726 N9726 N9727 Segment
X9727 N9727 N9728 Segment
X9728 N9728 N9729 Segment
X9729 N9729 N9730 Segment
X9730 N9730 N9731 Segment
X9731 N9731 N9732 Segment
X9732 N9732 N9733 Segment
X9733 N9733 N9734 Segment
X9734 N9734 N9735 Segment
X9735 N9735 N9736 Segment
X9736 N9736 N9737 Segment
X9737 N9737 N9738 Segment
X9738 N9738 N9739 Segment
X9739 N9739 N9740 Segment
X9740 N9740 N9741 Segment
X9741 N9741 N9742 Segment
X9742 N9742 N9743 Segment
X9743 N9743 N9744 Segment
X9744 N9744 N9745 Segment
X9745 N9745 N9746 Segment
X9746 N9746 N9747 Segment
X9747 N9747 N9748 Segment
X9748 N9748 N9749 Segment
X9749 N9749 N9750 Segment
X9750 N9750 N9751 Segment
X9751 N9751 N9752 Segment
X9752 N9752 N9753 Segment
X9753 N9753 N9754 Segment
X9754 N9754 N9755 Segment
X9755 N9755 N9756 Segment
X9756 N9756 N9757 Segment
X9757 N9757 N9758 Segment
X9758 N9758 N9759 Segment
X9759 N9759 N9760 Segment
X9760 N9760 N9761 Segment
X9761 N9761 N9762 Segment
X9762 N9762 N9763 Segment
X9763 N9763 N9764 Segment
X9764 N9764 N9765 Segment
X9765 N9765 N9766 Segment
X9766 N9766 N9767 Segment
X9767 N9767 N9768 Segment
X9768 N9768 N9769 Segment
X9769 N9769 N9770 Segment
X9770 N9770 N9771 Segment
X9771 N9771 N9772 Segment
X9772 N9772 N9773 Segment
X9773 N9773 N9774 Segment
X9774 N9774 N9775 Segment
X9775 N9775 N9776 Segment
X9776 N9776 N9777 Segment
X9777 N9777 N9778 Segment
X9778 N9778 N9779 Segment
X9779 N9779 N9780 Segment
X9780 N9780 N9781 Segment
X9781 N9781 N9782 Segment
X9782 N9782 N9783 Segment
X9783 N9783 N9784 Segment
X9784 N9784 N9785 Segment
X9785 N9785 N9786 Segment
X9786 N9786 N9787 Segment
X9787 N9787 N9788 Segment
X9788 N9788 N9789 Segment
X9789 N9789 N9790 Segment
X9790 N9790 N9791 Segment
X9791 N9791 N9792 Segment
X9792 N9792 N9793 Segment
X9793 N9793 N9794 Segment
X9794 N9794 N9795 Segment
X9795 N9795 N9796 Segment
X9796 N9796 N9797 Segment
X9797 N9797 N9798 Segment
X9798 N9798 N9799 Segment
X9799 N9799 N9800 Segment
X9800 N9800 N9801 Segment
X9801 N9801 N9802 Segment
X9802 N9802 N9803 Segment
X9803 N9803 N9804 Segment
X9804 N9804 N9805 Segment
X9805 N9805 N9806 Segment
X9806 N9806 N9807 Segment
X9807 N9807 N9808 Segment
X9808 N9808 N9809 Segment
X9809 N9809 N9810 Segment
X9810 N9810 N9811 Segment
X9811 N9811 N9812 Segment
X9812 N9812 N9813 Segment
X9813 N9813 N9814 Segment
X9814 N9814 N9815 Segment
X9815 N9815 N9816 Segment
X9816 N9816 N9817 Segment
X9817 N9817 N9818 Segment
X9818 N9818 N9819 Segment
X9819 N9819 N9820 Segment
X9820 N9820 N9821 Segment
X9821 N9821 N9822 Segment
X9822 N9822 N9823 Segment
X9823 N9823 N9824 Segment
X9824 N9824 N9825 Segment
X9825 N9825 N9826 Segment
X9826 N9826 N9827 Segment
X9827 N9827 N9828 Segment
X9828 N9828 N9829 Segment
X9829 N9829 N9830 Segment
X9830 N9830 N9831 Segment
X9831 N9831 N9832 Segment
X9832 N9832 N9833 Segment
X9833 N9833 N9834 Segment
X9834 N9834 N9835 Segment
X9835 N9835 N9836 Segment
X9836 N9836 N9837 Segment
X9837 N9837 N9838 Segment
X9838 N9838 N9839 Segment
X9839 N9839 N9840 Segment
X9840 N9840 N9841 Segment
X9841 N9841 N9842 Segment
X9842 N9842 N9843 Segment
X9843 N9843 N9844 Segment
X9844 N9844 N9845 Segment
X9845 N9845 N9846 Segment
X9846 N9846 N9847 Segment
X9847 N9847 N9848 Segment
X9848 N9848 N9849 Segment
X9849 N9849 N9850 Segment
X9850 N9850 N9851 Segment
X9851 N9851 N9852 Segment
X9852 N9852 N9853 Segment
X9853 N9853 N9854 Segment
X9854 N9854 N9855 Segment
X9855 N9855 N9856 Segment
X9856 N9856 N9857 Segment
X9857 N9857 N9858 Segment
X9858 N9858 N9859 Segment
X9859 N9859 N9860 Segment
X9860 N9860 N9861 Segment
X9861 N9861 N9862 Segment
X9862 N9862 N9863 Segment
X9863 N9863 N9864 Segment
X9864 N9864 N9865 Segment
X9865 N9865 N9866 Segment
X9866 N9866 N9867 Segment
X9867 N9867 N9868 Segment
X9868 N9868 N9869 Segment
X9869 N9869 N9870 Segment
X9870 N9870 N9871 Segment
X9871 N9871 N9872 Segment
X9872 N9872 N9873 Segment
X9873 N9873 N9874 Segment
X9874 N9874 N9875 Segment
X9875 N9875 N9876 Segment
X9876 N9876 N9877 Segment
X9877 N9877 N9878 Segment
X9878 N9878 N9879 Segment
X9879 N9879 N9880 Segment
X9880 N9880 N9881 Segment
X9881 N9881 N9882 Segment
X9882 N9882 N9883 Segment
X9883 N9883 N9884 Segment
X9884 N9884 N9885 Segment
X9885 N9885 N9886 Segment
X9886 N9886 N9887 Segment
X9887 N9887 N9888 Segment
X9888 N9888 N9889 Segment
X9889 N9889 N9890 Segment
X9890 N9890 N9891 Segment
X9891 N9891 N9892 Segment
X9892 N9892 N9893 Segment
X9893 N9893 N9894 Segment
X9894 N9894 N9895 Segment
X9895 N9895 N9896 Segment
X9896 N9896 N9897 Segment
X9897 N9897 N9898 Segment
X9898 N9898 N9899 Segment
X9899 N9899 N9900 Segment
X9900 N9900 N9901 Segment
X9901 N9901 N9902 Segment
X9902 N9902 N9903 Segment
X9903 N9903 N9904 Segment
X9904 N9904 N9905 Segment
X9905 N9905 N9906 Segment
X9906 N9906 N9907 Segment
X9907 N9907 N9908 Segment
X9908 N9908 N9909 Segment
X9909 N9909 N9910 Segment
X9910 N9910 N9911 Segment
X9911 N9911 N9912 Segment
X9912 N9912 N9913 Segment
X9913 N9913 N9914 Segment
X9914 N9914 N9915 Segment
X9915 N9915 N9916 Segment
X9916 N9916 N9917 Segment
X9917 N9917 N9918 Segment
X9918 N9918 N9919 Segment
X9919 N9919 N9920 Segment
X9920 N9920 N9921 Segment
X9921 N9921 N9922 Segment
X9922 N9922 N9923 Segment
X9923 N9923 N9924 Segment
X9924 N9924 N9925 Segment
X9925 N9925 N9926 Segment
X9926 N9926 N9927 Segment
X9927 N9927 N9928 Segment
X9928 N9928 N9929 Segment
X9929 N9929 N9930 Segment
X9930 N9930 N9931 Segment
X9931 N9931 N9932 Segment
X9932 N9932 N9933 Segment
X9933 N9933 N9934 Segment
X9934 N9934 N9935 Segment
X9935 N9935 N9936 Segment
X9936 N9936 N9937 Segment
X9937 N9937 N9938 Segment
X9938 N9938 N9939 Segment
X9939 N9939 N9940 Segment
X9940 N9940 N9941 Segment
X9941 N9941 N9942 Segment
X9942 N9942 N9943 Segment
X9943 N9943 N9944 Segment
X9944 N9944 N9945 Segment
X9945 N9945 N9946 Segment
X9946 N9946 N9947 Segment
X9947 N9947 N9948 Segment
X9948 N9948 N9949 Segment
X9949 N9949 N9950 Segment
X9950 N9950 N9951 Segment
X9951 N9951 N9952 Segment
X9952 N9952 N9953 Segment
X9953 N9953 N9954 Segment
X9954 N9954 N9955 Segment
X9955 N9955 N9956 Segment
X9956 N9956 N9957 Segment
X9957 N9957 N9958 Segment
X9958 N9958 N9959 Segment
X9959 N9959 N9960 Segment
X9960 N9960 N9961 Segment
X9961 N9961 N9962 Segment
X9962 N9962 N9963 Segment
X9963 N9963 N9964 Segment
X9964 N9964 N9965 Segment
X9965 N9965 N9966 Segment
X9966 N9966 N9967 Segment
X9967 N9967 N9968 Segment
X9968 N9968 N9969 Segment
X9969 N9969 N9970 Segment
X9970 N9970 N9971 Segment
X9971 N9971 N9972 Segment
X9972 N9972 N9973 Segment
X9973 N9973 N9974 Segment
X9974 N9974 N9975 Segment
X9975 N9975 N9976 Segment
X9976 N9976 N9977 Segment
X9977 N9977 N9978 Segment
X9978 N9978 N9979 Segment
X9979 N9979 N9980 Segment
X9980 N9980 N9981 Segment
X9981 N9981 N9982 Segment
X9982 N9982 N9983 Segment
X9983 N9983 N9984 Segment
X9984 N9984 N9985 Segment
X9985 N9985 N9986 Segment
X9986 N9986 N9987 Segment
X9987 N9987 N9988 Segment
X9988 N9988 N9989 Segment
X9989 N9989 N9990 Segment
X9990 N9990 N9991 Segment
X9991 N9991 N9992 Segment
X9992 N9992 N9993 Segment
X9993 N9993 N9994 Segment
X9994 N9994 N9995 Segment
X9995 N9995 N9996 Segment
X9996 N9996 N9997 Segment
X9997 N9997 N9998 Segment
X9998 N9998 N9999 Segment
X9999 N9999 N10000 Segment
X10000 N10000 N10001 Segment
X10001 N10001 N10002 Segment
X10002 N10002 N10003 Segment
X10003 N10003 N10004 Segment
X10004 N10004 N10005 Segment
X10005 N10005 N10006 Segment
X10006 N10006 N10007 Segment
X10007 N10007 N10008 Segment
X10008 N10008 N10009 Segment
X10009 N10009 N10010 Segment
X10010 N10010 N10011 Segment
X10011 N10011 N10012 Segment
X10012 N10012 N10013 Segment
X10013 N10013 N10014 Segment
X10014 N10014 N10015 Segment
X10015 N10015 N10016 Segment
X10016 N10016 N10017 Segment
X10017 N10017 N10018 Segment
X10018 N10018 N10019 Segment
X10019 N10019 N10020 Segment
X10020 N10020 N10021 Segment
X10021 N10021 N10022 Segment
X10022 N10022 N10023 Segment
X10023 N10023 N10024 Segment
X10024 N10024 N10025 Segment
X10025 N10025 N10026 Segment
X10026 N10026 N10027 Segment
X10027 N10027 N10028 Segment
X10028 N10028 N10029 Segment
X10029 N10029 N10030 Segment
X10030 N10030 N10031 Segment
X10031 N10031 N10032 Segment
X10032 N10032 N10033 Segment
X10033 N10033 N10034 Segment
X10034 N10034 N10035 Segment
X10035 N10035 N10036 Segment
X10036 N10036 N10037 Segment
X10037 N10037 N10038 Segment
X10038 N10038 N10039 Segment
X10039 N10039 N10040 Segment
X10040 N10040 N10041 Segment
X10041 N10041 N10042 Segment
X10042 N10042 N10043 Segment
X10043 N10043 N10044 Segment
X10044 N10044 N10045 Segment
X10045 N10045 N10046 Segment
X10046 N10046 N10047 Segment
X10047 N10047 N10048 Segment
X10048 N10048 N10049 Segment
X10049 N10049 N10050 Segment
X10050 N10050 N10051 Segment
X10051 N10051 N10052 Segment
X10052 N10052 N10053 Segment
X10053 N10053 N10054 Segment
X10054 N10054 N10055 Segment
X10055 N10055 N10056 Segment
X10056 N10056 N10057 Segment
X10057 N10057 N10058 Segment
X10058 N10058 N10059 Segment
X10059 N10059 N10060 Segment
X10060 N10060 N10061 Segment
X10061 N10061 N10062 Segment
X10062 N10062 N10063 Segment
X10063 N10063 N10064 Segment
X10064 N10064 N10065 Segment
X10065 N10065 N10066 Segment
X10066 N10066 N10067 Segment
X10067 N10067 N10068 Segment
X10068 N10068 N10069 Segment
X10069 N10069 N10070 Segment
X10070 N10070 N10071 Segment
X10071 N10071 N10072 Segment
X10072 N10072 N10073 Segment
X10073 N10073 N10074 Segment
X10074 N10074 N10075 Segment
X10075 N10075 N10076 Segment
X10076 N10076 N10077 Segment
X10077 N10077 N10078 Segment
X10078 N10078 N10079 Segment
X10079 N10079 N10080 Segment
X10080 N10080 N10081 Segment
X10081 N10081 N10082 Segment
X10082 N10082 N10083 Segment
X10083 N10083 N10084 Segment
X10084 N10084 N10085 Segment
X10085 N10085 N10086 Segment
X10086 N10086 N10087 Segment
X10087 N10087 N10088 Segment
X10088 N10088 N10089 Segment
X10089 N10089 N10090 Segment
X10090 N10090 N10091 Segment
X10091 N10091 N10092 Segment
X10092 N10092 N10093 Segment
X10093 N10093 N10094 Segment
X10094 N10094 N10095 Segment
X10095 N10095 N10096 Segment
X10096 N10096 N10097 Segment
X10097 N10097 N10098 Segment
X10098 N10098 N10099 Segment
X10099 N10099 N10100 Segment
X10100 N10100 N10101 Segment
X10101 N10101 N10102 Segment
X10102 N10102 N10103 Segment
X10103 N10103 N10104 Segment
X10104 N10104 N10105 Segment
X10105 N10105 N10106 Segment
X10106 N10106 N10107 Segment
X10107 N10107 N10108 Segment
X10108 N10108 N10109 Segment
X10109 N10109 N10110 Segment
X10110 N10110 N10111 Segment
X10111 N10111 N10112 Segment
X10112 N10112 N10113 Segment
X10113 N10113 N10114 Segment
X10114 N10114 N10115 Segment
X10115 N10115 N10116 Segment
X10116 N10116 N10117 Segment
X10117 N10117 N10118 Segment
X10118 N10118 N10119 Segment
X10119 N10119 N10120 Segment
X10120 N10120 N10121 Segment
X10121 N10121 N10122 Segment
X10122 N10122 N10123 Segment
X10123 N10123 N10124 Segment
X10124 N10124 N10125 Segment
X10125 N10125 N10126 Segment
X10126 N10126 N10127 Segment
X10127 N10127 N10128 Segment
X10128 N10128 N10129 Segment
X10129 N10129 N10130 Segment
X10130 N10130 N10131 Segment
X10131 N10131 N10132 Segment
X10132 N10132 N10133 Segment
X10133 N10133 N10134 Segment
X10134 N10134 N10135 Segment
X10135 N10135 N10136 Segment
X10136 N10136 N10137 Segment
X10137 N10137 N10138 Segment
X10138 N10138 N10139 Segment
X10139 N10139 N10140 Segment
X10140 N10140 N10141 Segment
X10141 N10141 N10142 Segment
X10142 N10142 N10143 Segment
X10143 N10143 N10144 Segment
X10144 N10144 N10145 Segment
X10145 N10145 N10146 Segment
X10146 N10146 N10147 Segment
X10147 N10147 N10148 Segment
X10148 N10148 N10149 Segment
X10149 N10149 N10150 Segment
X10150 N10150 N10151 Segment
X10151 N10151 N10152 Segment
X10152 N10152 N10153 Segment
X10153 N10153 N10154 Segment
X10154 N10154 N10155 Segment
X10155 N10155 N10156 Segment
X10156 N10156 N10157 Segment
X10157 N10157 N10158 Segment
X10158 N10158 N10159 Segment
X10159 N10159 N10160 Segment
X10160 N10160 N10161 Segment
X10161 N10161 N10162 Segment
X10162 N10162 N10163 Segment
X10163 N10163 N10164 Segment
X10164 N10164 N10165 Segment
X10165 N10165 N10166 Segment
X10166 N10166 N10167 Segment
X10167 N10167 N10168 Segment
X10168 N10168 N10169 Segment
X10169 N10169 N10170 Segment
X10170 N10170 N10171 Segment
X10171 N10171 N10172 Segment
X10172 N10172 N10173 Segment
X10173 N10173 N10174 Segment
X10174 N10174 N10175 Segment
X10175 N10175 N10176 Segment
X10176 N10176 N10177 Segment
X10177 N10177 N10178 Segment
X10178 N10178 N10179 Segment
X10179 N10179 N10180 Segment
X10180 N10180 N10181 Segment
X10181 N10181 N10182 Segment
X10182 N10182 N10183 Segment
X10183 N10183 N10184 Segment
X10184 N10184 N10185 Segment
X10185 N10185 N10186 Segment
X10186 N10186 N10187 Segment
X10187 N10187 N10188 Segment
X10188 N10188 N10189 Segment
X10189 N10189 N10190 Segment
X10190 N10190 N10191 Segment
X10191 N10191 N10192 Segment
X10192 N10192 N10193 Segment
X10193 N10193 N10194 Segment
X10194 N10194 N10195 Segment
X10195 N10195 N10196 Segment
X10196 N10196 N10197 Segment
X10197 N10197 N10198 Segment
X10198 N10198 N10199 Segment
X10199 N10199 N10200 Segment
X10200 N10200 N10201 Segment
X10201 N10201 N10202 Segment
X10202 N10202 N10203 Segment
X10203 N10203 N10204 Segment
X10204 N10204 N10205 Segment
X10205 N10205 N10206 Segment
X10206 N10206 N10207 Segment
X10207 N10207 N10208 Segment
X10208 N10208 N10209 Segment
X10209 N10209 N10210 Segment
X10210 N10210 N10211 Segment
X10211 N10211 N10212 Segment
X10212 N10212 N10213 Segment
X10213 N10213 N10214 Segment
X10214 N10214 N10215 Segment
X10215 N10215 N10216 Segment
X10216 N10216 N10217 Segment
X10217 N10217 N10218 Segment
X10218 N10218 N10219 Segment
X10219 N10219 N10220 Segment
X10220 N10220 N10221 Segment
X10221 N10221 N10222 Segment
X10222 N10222 N10223 Segment
X10223 N10223 N10224 Segment
X10224 N10224 N10225 Segment
X10225 N10225 N10226 Segment
X10226 N10226 N10227 Segment
X10227 N10227 N10228 Segment
X10228 N10228 N10229 Segment
X10229 N10229 N10230 Segment
X10230 N10230 N10231 Segment
X10231 N10231 N10232 Segment
X10232 N10232 N10233 Segment
X10233 N10233 N10234 Segment
X10234 N10234 N10235 Segment
X10235 N10235 N10236 Segment
X10236 N10236 N10237 Segment
X10237 N10237 N10238 Segment
X10238 N10238 N10239 Segment
X10239 N10239 N10240 Segment
X10240 N10240 N10241 Segment
X10241 N10241 N10242 Segment
X10242 N10242 N10243 Segment
X10243 N10243 N10244 Segment
X10244 N10244 N10245 Segment
X10245 N10245 N10246 Segment
X10246 N10246 N10247 Segment
X10247 N10247 N10248 Segment
X10248 N10248 N10249 Segment
X10249 N10249 N10250 Segment
X10250 N10250 N10251 Segment
X10251 N10251 N10252 Segment
X10252 N10252 N10253 Segment
X10253 N10253 N10254 Segment
X10254 N10254 N10255 Segment
X10255 N10255 N10256 Segment
X10256 N10256 N10257 Segment
X10257 N10257 N10258 Segment
X10258 N10258 N10259 Segment
X10259 N10259 N10260 Segment
X10260 N10260 N10261 Segment
X10261 N10261 N10262 Segment
X10262 N10262 N10263 Segment
X10263 N10263 N10264 Segment
X10264 N10264 N10265 Segment
X10265 N10265 N10266 Segment
X10266 N10266 N10267 Segment
X10267 N10267 N10268 Segment
X10268 N10268 N10269 Segment
X10269 N10269 N10270 Segment
X10270 N10270 N10271 Segment
X10271 N10271 N10272 Segment
X10272 N10272 N10273 Segment
X10273 N10273 N10274 Segment
X10274 N10274 N10275 Segment
X10275 N10275 N10276 Segment
X10276 N10276 N10277 Segment
X10277 N10277 N10278 Segment
X10278 N10278 N10279 Segment
X10279 N10279 N10280 Segment
X10280 N10280 N10281 Segment
X10281 N10281 N10282 Segment
X10282 N10282 N10283 Segment
X10283 N10283 N10284 Segment
X10284 N10284 N10285 Segment
X10285 N10285 N10286 Segment
X10286 N10286 N10287 Segment
X10287 N10287 N10288 Segment
X10288 N10288 N10289 Segment
X10289 N10289 N10290 Segment
X10290 N10290 N10291 Segment
X10291 N10291 N10292 Segment
X10292 N10292 N10293 Segment
X10293 N10293 N10294 Segment
X10294 N10294 N10295 Segment
X10295 N10295 N10296 Segment
X10296 N10296 N10297 Segment
X10297 N10297 N10298 Segment
X10298 N10298 N10299 Segment
X10299 N10299 N10300 Segment
X10300 N10300 N10301 Segment
X10301 N10301 N10302 Segment
X10302 N10302 N10303 Segment
X10303 N10303 N10304 Segment
X10304 N10304 N10305 Segment
X10305 N10305 N10306 Segment
X10306 N10306 N10307 Segment
X10307 N10307 N10308 Segment
X10308 N10308 N10309 Segment
X10309 N10309 N10310 Segment
X10310 N10310 N10311 Segment
X10311 N10311 N10312 Segment
X10312 N10312 N10313 Segment
X10313 N10313 N10314 Segment
X10314 N10314 N10315 Segment
X10315 N10315 N10316 Segment
X10316 N10316 N10317 Segment
X10317 N10317 N10318 Segment
X10318 N10318 N10319 Segment
X10319 N10319 N10320 Segment
X10320 N10320 N10321 Segment
X10321 N10321 N10322 Segment
X10322 N10322 N10323 Segment
X10323 N10323 N10324 Segment
X10324 N10324 N10325 Segment
X10325 N10325 N10326 Segment
X10326 N10326 N10327 Segment
X10327 N10327 N10328 Segment
X10328 N10328 N10329 Segment
X10329 N10329 N10330 Segment
X10330 N10330 N10331 Segment
X10331 N10331 N10332 Segment
X10332 N10332 N10333 Segment
X10333 N10333 N10334 Segment
X10334 N10334 N10335 Segment
X10335 N10335 N10336 Segment
X10336 N10336 N10337 Segment
X10337 N10337 N10338 Segment
X10338 N10338 N10339 Segment
X10339 N10339 N10340 Segment
X10340 N10340 N10341 Segment
X10341 N10341 N10342 Segment
X10342 N10342 N10343 Segment
X10343 N10343 N10344 Segment
X10344 N10344 N10345 Segment
X10345 N10345 N10346 Segment
X10346 N10346 N10347 Segment
X10347 N10347 N10348 Segment
X10348 N10348 N10349 Segment
X10349 N10349 N10350 Segment
X10350 N10350 N10351 Segment
X10351 N10351 N10352 Segment
X10352 N10352 N10353 Segment
X10353 N10353 N10354 Segment
X10354 N10354 N10355 Segment
X10355 N10355 N10356 Segment
X10356 N10356 N10357 Segment
X10357 N10357 N10358 Segment
X10358 N10358 N10359 Segment
X10359 N10359 N10360 Segment
X10360 N10360 N10361 Segment
X10361 N10361 N10362 Segment
X10362 N10362 N10363 Segment
X10363 N10363 N10364 Segment
X10364 N10364 N10365 Segment
X10365 N10365 N10366 Segment
X10366 N10366 N10367 Segment
X10367 N10367 N10368 Segment
X10368 N10368 N10369 Segment
X10369 N10369 N10370 Segment
X10370 N10370 N10371 Segment
X10371 N10371 N10372 Segment
X10372 N10372 N10373 Segment
X10373 N10373 N10374 Segment
X10374 N10374 N10375 Segment
X10375 N10375 N10376 Segment
X10376 N10376 N10377 Segment
X10377 N10377 N10378 Segment
X10378 N10378 N10379 Segment
X10379 N10379 N10380 Segment
X10380 N10380 N10381 Segment
X10381 N10381 N10382 Segment
X10382 N10382 N10383 Segment
X10383 N10383 N10384 Segment
X10384 N10384 N10385 Segment
X10385 N10385 N10386 Segment
X10386 N10386 N10387 Segment
X10387 N10387 N10388 Segment
X10388 N10388 N10389 Segment
X10389 N10389 N10390 Segment
X10390 N10390 N10391 Segment
X10391 N10391 N10392 Segment
X10392 N10392 N10393 Segment
X10393 N10393 N10394 Segment
X10394 N10394 N10395 Segment
X10395 N10395 N10396 Segment
X10396 N10396 N10397 Segment
X10397 N10397 N10398 Segment
X10398 N10398 N10399 Segment
X10399 N10399 N10400 Segment
X10400 N10400 N10401 Segment
X10401 N10401 N10402 Segment
X10402 N10402 N10403 Segment
X10403 N10403 N10404 Segment
X10404 N10404 N10405 Segment
X10405 N10405 N10406 Segment
X10406 N10406 N10407 Segment
X10407 N10407 N10408 Segment
X10408 N10408 N10409 Segment
X10409 N10409 N10410 Segment
X10410 N10410 N10411 Segment
X10411 N10411 N10412 Segment
X10412 N10412 N10413 Segment
X10413 N10413 N10414 Segment
X10414 N10414 N10415 Segment
X10415 N10415 N10416 Segment
X10416 N10416 N10417 Segment
X10417 N10417 N10418 Segment
X10418 N10418 N10419 Segment
X10419 N10419 N10420 Segment
X10420 N10420 N10421 Segment
X10421 N10421 N10422 Segment
X10422 N10422 N10423 Segment
X10423 N10423 N10424 Segment
X10424 N10424 N10425 Segment
X10425 N10425 N10426 Segment
X10426 N10426 N10427 Segment
X10427 N10427 N10428 Segment
X10428 N10428 N10429 Segment
X10429 N10429 N10430 Segment
X10430 N10430 N10431 Segment
X10431 N10431 N10432 Segment
X10432 N10432 N10433 Segment
X10433 N10433 N10434 Segment
X10434 N10434 N10435 Segment
X10435 N10435 N10436 Segment
X10436 N10436 N10437 Segment
X10437 N10437 N10438 Segment
X10438 N10438 N10439 Segment
X10439 N10439 N10440 Segment
X10440 N10440 N10441 Segment
X10441 N10441 N10442 Segment
X10442 N10442 N10443 Segment
X10443 N10443 N10444 Segment
X10444 N10444 N10445 Segment
X10445 N10445 N10446 Segment
X10446 N10446 N10447 Segment
X10447 N10447 N10448 Segment
X10448 N10448 N10449 Segment
X10449 N10449 N10450 Segment
X10450 N10450 N10451 Segment
X10451 N10451 N10452 Segment
X10452 N10452 N10453 Segment
X10453 N10453 N10454 Segment
X10454 N10454 N10455 Segment
X10455 N10455 N10456 Segment
X10456 N10456 N10457 Segment
X10457 N10457 N10458 Segment
X10458 N10458 N10459 Segment
X10459 N10459 N10460 Segment
X10460 N10460 N10461 Segment
X10461 N10461 N10462 Segment
X10462 N10462 N10463 Segment
X10463 N10463 N10464 Segment
X10464 N10464 N10465 Segment
X10465 N10465 N10466 Segment
X10466 N10466 N10467 Segment
X10467 N10467 N10468 Segment
X10468 N10468 N10469 Segment
X10469 N10469 N10470 Segment
X10470 N10470 N10471 Segment
X10471 N10471 N10472 Segment
X10472 N10472 N10473 Segment
X10473 N10473 N10474 Segment
X10474 N10474 N10475 Segment
X10475 N10475 N10476 Segment
X10476 N10476 N10477 Segment
X10477 N10477 N10478 Segment
X10478 N10478 N10479 Segment
X10479 N10479 N10480 Segment
X10480 N10480 N10481 Segment
X10481 N10481 N10482 Segment
X10482 N10482 N10483 Segment
X10483 N10483 N10484 Segment
X10484 N10484 N10485 Segment
X10485 N10485 N10486 Segment
X10486 N10486 N10487 Segment
X10487 N10487 N10488 Segment
X10488 N10488 N10489 Segment
X10489 N10489 N10490 Segment
X10490 N10490 N10491 Segment
X10491 N10491 N10492 Segment
X10492 N10492 N10493 Segment
X10493 N10493 N10494 Segment
X10494 N10494 N10495 Segment
X10495 N10495 N10496 Segment
X10496 N10496 N10497 Segment
X10497 N10497 N10498 Segment
X10498 N10498 N10499 Segment
X10499 N10499 N10500 Segment
X10500 N10500 N10501 Segment
X10501 N10501 N10502 Segment
X10502 N10502 N10503 Segment
X10503 N10503 N10504 Segment
X10504 N10504 N10505 Segment
X10505 N10505 N10506 Segment
X10506 N10506 N10507 Segment
X10507 N10507 N10508 Segment
X10508 N10508 N10509 Segment
X10509 N10509 N10510 Segment
X10510 N10510 N10511 Segment
X10511 N10511 N10512 Segment
X10512 N10512 N10513 Segment
X10513 N10513 N10514 Segment
X10514 N10514 N10515 Segment
X10515 N10515 N10516 Segment
X10516 N10516 N10517 Segment
X10517 N10517 N10518 Segment
X10518 N10518 N10519 Segment
X10519 N10519 N10520 Segment
X10520 N10520 N10521 Segment
X10521 N10521 N10522 Segment
X10522 N10522 N10523 Segment
X10523 N10523 N10524 Segment
X10524 N10524 N10525 Segment
X10525 N10525 N10526 Segment
X10526 N10526 N10527 Segment
X10527 N10527 N10528 Segment
X10528 N10528 N10529 Segment
X10529 N10529 N10530 Segment
X10530 N10530 N10531 Segment
X10531 N10531 N10532 Segment
X10532 N10532 N10533 Segment
X10533 N10533 N10534 Segment
X10534 N10534 N10535 Segment
X10535 N10535 N10536 Segment
X10536 N10536 N10537 Segment
X10537 N10537 N10538 Segment
X10538 N10538 N10539 Segment
X10539 N10539 N10540 Segment
X10540 N10540 N10541 Segment
X10541 N10541 N10542 Segment
X10542 N10542 N10543 Segment
X10543 N10543 N10544 Segment
X10544 N10544 N10545 Segment
X10545 N10545 N10546 Segment
X10546 N10546 N10547 Segment
X10547 N10547 N10548 Segment
X10548 N10548 N10549 Segment
X10549 N10549 N10550 Segment
X10550 N10550 N10551 Segment
X10551 N10551 N10552 Segment
X10552 N10552 N10553 Segment
X10553 N10553 N10554 Segment
X10554 N10554 N10555 Segment
X10555 N10555 N10556 Segment
X10556 N10556 N10557 Segment
X10557 N10557 N10558 Segment
X10558 N10558 N10559 Segment
X10559 N10559 N10560 Segment
X10560 N10560 N10561 Segment
X10561 N10561 N10562 Segment
X10562 N10562 N10563 Segment
X10563 N10563 N10564 Segment
X10564 N10564 N10565 Segment
X10565 N10565 N10566 Segment
X10566 N10566 N10567 Segment
X10567 N10567 N10568 Segment
X10568 N10568 N10569 Segment
X10569 N10569 N10570 Segment
X10570 N10570 N10571 Segment
X10571 N10571 N10572 Segment
X10572 N10572 N10573 Segment
X10573 N10573 N10574 Segment
X10574 N10574 N10575 Segment
X10575 N10575 N10576 Segment
X10576 N10576 N10577 Segment
X10577 N10577 N10578 Segment
X10578 N10578 N10579 Segment
X10579 N10579 N10580 Segment
X10580 N10580 N10581 Segment
X10581 N10581 N10582 Segment
X10582 N10582 N10583 Segment
X10583 N10583 N10584 Segment
X10584 N10584 N10585 Segment
X10585 N10585 N10586 Segment
X10586 N10586 N10587 Segment
X10587 N10587 N10588 Segment
X10588 N10588 N10589 Segment
X10589 N10589 N10590 Segment
X10590 N10590 N10591 Segment
X10591 N10591 N10592 Segment
X10592 N10592 N10593 Segment
X10593 N10593 N10594 Segment
X10594 N10594 N10595 Segment
X10595 N10595 N10596 Segment
X10596 N10596 N10597 Segment
X10597 N10597 N10598 Segment
X10598 N10598 N10599 Segment
X10599 N10599 N10600 Segment
X10600 N10600 N10601 Segment
X10601 N10601 N10602 Segment
X10602 N10602 N10603 Segment
X10603 N10603 N10604 Segment
X10604 N10604 N10605 Segment
X10605 N10605 N10606 Segment
X10606 N10606 N10607 Segment
X10607 N10607 N10608 Segment
X10608 N10608 N10609 Segment
X10609 N10609 N10610 Segment
X10610 N10610 N10611 Segment
X10611 N10611 N10612 Segment
X10612 N10612 N10613 Segment
X10613 N10613 N10614 Segment
X10614 N10614 N10615 Segment
X10615 N10615 N10616 Segment
X10616 N10616 N10617 Segment
X10617 N10617 N10618 Segment
X10618 N10618 N10619 Segment
X10619 N10619 N10620 Segment
X10620 N10620 N10621 Segment
X10621 N10621 N10622 Segment
X10622 N10622 N10623 Segment
X10623 N10623 N10624 Segment
X10624 N10624 N10625 Segment
X10625 N10625 N10626 Segment
X10626 N10626 N10627 Segment
X10627 N10627 N10628 Segment
X10628 N10628 N10629 Segment
X10629 N10629 N10630 Segment
X10630 N10630 N10631 Segment
X10631 N10631 N10632 Segment
X10632 N10632 N10633 Segment
X10633 N10633 N10634 Segment
X10634 N10634 N10635 Segment
X10635 N10635 N10636 Segment
X10636 N10636 N10637 Segment
X10637 N10637 N10638 Segment
X10638 N10638 N10639 Segment
X10639 N10639 N10640 Segment
X10640 N10640 N10641 Segment
X10641 N10641 N10642 Segment
X10642 N10642 N10643 Segment
X10643 N10643 N10644 Segment
X10644 N10644 N10645 Segment
X10645 N10645 N10646 Segment
X10646 N10646 N10647 Segment
X10647 N10647 N10648 Segment
X10648 N10648 N10649 Segment
X10649 N10649 N10650 Segment
X10650 N10650 N10651 Segment
X10651 N10651 N10652 Segment
X10652 N10652 N10653 Segment
X10653 N10653 N10654 Segment
X10654 N10654 N10655 Segment
X10655 N10655 N10656 Segment
X10656 N10656 N10657 Segment
X10657 N10657 N10658 Segment
X10658 N10658 N10659 Segment
X10659 N10659 N10660 Segment
X10660 N10660 N10661 Segment
X10661 N10661 N10662 Segment
X10662 N10662 N10663 Segment
X10663 N10663 N10664 Segment
X10664 N10664 N10665 Segment
X10665 N10665 N10666 Segment
X10666 N10666 N10667 Segment
X10667 N10667 N10668 Segment
X10668 N10668 N10669 Segment
X10669 N10669 N10670 Segment
X10670 N10670 N10671 Segment
X10671 N10671 N10672 Segment
X10672 N10672 N10673 Segment
X10673 N10673 N10674 Segment
X10674 N10674 N10675 Segment
X10675 N10675 N10676 Segment
X10676 N10676 N10677 Segment
X10677 N10677 N10678 Segment
X10678 N10678 N10679 Segment
X10679 N10679 N10680 Segment
X10680 N10680 N10681 Segment
X10681 N10681 N10682 Segment
X10682 N10682 N10683 Segment
X10683 N10683 N10684 Segment
X10684 N10684 N10685 Segment
X10685 N10685 N10686 Segment
X10686 N10686 N10687 Segment
X10687 N10687 N10688 Segment
X10688 N10688 N10689 Segment
X10689 N10689 N10690 Segment
X10690 N10690 N10691 Segment
X10691 N10691 N10692 Segment
X10692 N10692 N10693 Segment
X10693 N10693 N10694 Segment
X10694 N10694 N10695 Segment
X10695 N10695 N10696 Segment
X10696 N10696 N10697 Segment
X10697 N10697 N10698 Segment
X10698 N10698 N10699 Segment
X10699 N10699 N10700 Segment
X10700 N10700 N10701 Segment
X10701 N10701 N10702 Segment
X10702 N10702 N10703 Segment
X10703 N10703 N10704 Segment
X10704 N10704 N10705 Segment
X10705 N10705 N10706 Segment
X10706 N10706 N10707 Segment
X10707 N10707 N10708 Segment
X10708 N10708 N10709 Segment
X10709 N10709 N10710 Segment
X10710 N10710 N10711 Segment
X10711 N10711 N10712 Segment
X10712 N10712 N10713 Segment
X10713 N10713 N10714 Segment
X10714 N10714 N10715 Segment
X10715 N10715 N10716 Segment
X10716 N10716 N10717 Segment
X10717 N10717 N10718 Segment
X10718 N10718 N10719 Segment
X10719 N10719 N10720 Segment
X10720 N10720 N10721 Segment
X10721 N10721 N10722 Segment
X10722 N10722 N10723 Segment
X10723 N10723 N10724 Segment
X10724 N10724 N10725 Segment
X10725 N10725 N10726 Segment
X10726 N10726 N10727 Segment
X10727 N10727 N10728 Segment
X10728 N10728 N10729 Segment
X10729 N10729 N10730 Segment
X10730 N10730 N10731 Segment
X10731 N10731 N10732 Segment
X10732 N10732 N10733 Segment
X10733 N10733 N10734 Segment
X10734 N10734 N10735 Segment
X10735 N10735 N10736 Segment
X10736 N10736 N10737 Segment
X10737 N10737 N10738 Segment
X10738 N10738 N10739 Segment
X10739 N10739 N10740 Segment
X10740 N10740 N10741 Segment
X10741 N10741 N10742 Segment
X10742 N10742 N10743 Segment
X10743 N10743 N10744 Segment
X10744 N10744 N10745 Segment
X10745 N10745 N10746 Segment
X10746 N10746 N10747 Segment
X10747 N10747 N10748 Segment
X10748 N10748 N10749 Segment
X10749 N10749 N10750 Segment
X10750 N10750 N10751 Segment
X10751 N10751 N10752 Segment
X10752 N10752 N10753 Segment
X10753 N10753 N10754 Segment
X10754 N10754 N10755 Segment
X10755 N10755 N10756 Segment
X10756 N10756 N10757 Segment
X10757 N10757 N10758 Segment
X10758 N10758 N10759 Segment
X10759 N10759 N10760 Segment
X10760 N10760 N10761 Segment
X10761 N10761 N10762 Segment
X10762 N10762 N10763 Segment
X10763 N10763 N10764 Segment
X10764 N10764 N10765 Segment
X10765 N10765 N10766 Segment
X10766 N10766 N10767 Segment
X10767 N10767 N10768 Segment
X10768 N10768 N10769 Segment
X10769 N10769 N10770 Segment
X10770 N10770 N10771 Segment
X10771 N10771 N10772 Segment
X10772 N10772 N10773 Segment
X10773 N10773 N10774 Segment
X10774 N10774 N10775 Segment
X10775 N10775 N10776 Segment
X10776 N10776 N10777 Segment
X10777 N10777 N10778 Segment
X10778 N10778 N10779 Segment
X10779 N10779 N10780 Segment
X10780 N10780 N10781 Segment
X10781 N10781 N10782 Segment
X10782 N10782 N10783 Segment
X10783 N10783 N10784 Segment
X10784 N10784 N10785 Segment
X10785 N10785 N10786 Segment
X10786 N10786 N10787 Segment
X10787 N10787 N10788 Segment
X10788 N10788 N10789 Segment
X10789 N10789 N10790 Segment
X10790 N10790 N10791 Segment
X10791 N10791 N10792 Segment
X10792 N10792 N10793 Segment
X10793 N10793 N10794 Segment
X10794 N10794 N10795 Segment
X10795 N10795 N10796 Segment
X10796 N10796 N10797 Segment
X10797 N10797 N10798 Segment
X10798 N10798 N10799 Segment
X10799 N10799 N10800 Segment
X10800 N10800 N10801 Segment
X10801 N10801 N10802 Segment
X10802 N10802 N10803 Segment
X10803 N10803 N10804 Segment
X10804 N10804 N10805 Segment
X10805 N10805 N10806 Segment
X10806 N10806 N10807 Segment
X10807 N10807 N10808 Segment
X10808 N10808 N10809 Segment
X10809 N10809 N10810 Segment
X10810 N10810 N10811 Segment
X10811 N10811 N10812 Segment
X10812 N10812 N10813 Segment
X10813 N10813 N10814 Segment
X10814 N10814 N10815 Segment
X10815 N10815 N10816 Segment
X10816 N10816 N10817 Segment
X10817 N10817 N10818 Segment
X10818 N10818 N10819 Segment
X10819 N10819 N10820 Segment
X10820 N10820 N10821 Segment
X10821 N10821 N10822 Segment
X10822 N10822 N10823 Segment
X10823 N10823 N10824 Segment
X10824 N10824 N10825 Segment
X10825 N10825 N10826 Segment
X10826 N10826 N10827 Segment
X10827 N10827 N10828 Segment
X10828 N10828 N10829 Segment
X10829 N10829 N10830 Segment
X10830 N10830 N10831 Segment
X10831 N10831 N10832 Segment
X10832 N10832 N10833 Segment
X10833 N10833 N10834 Segment
X10834 N10834 N10835 Segment
X10835 N10835 N10836 Segment
X10836 N10836 N10837 Segment
X10837 N10837 N10838 Segment
X10838 N10838 N10839 Segment
X10839 N10839 N10840 Segment
X10840 N10840 N10841 Segment
X10841 N10841 N10842 Segment
X10842 N10842 N10843 Segment
X10843 N10843 N10844 Segment
X10844 N10844 N10845 Segment
X10845 N10845 N10846 Segment
X10846 N10846 N10847 Segment
X10847 N10847 N10848 Segment
X10848 N10848 N10849 Segment
X10849 N10849 N10850 Segment
X10850 N10850 N10851 Segment
X10851 N10851 N10852 Segment
X10852 N10852 N10853 Segment
X10853 N10853 N10854 Segment
X10854 N10854 N10855 Segment
X10855 N10855 N10856 Segment
X10856 N10856 N10857 Segment
X10857 N10857 N10858 Segment
X10858 N10858 N10859 Segment
X10859 N10859 N10860 Segment
X10860 N10860 N10861 Segment
X10861 N10861 N10862 Segment
X10862 N10862 N10863 Segment
X10863 N10863 N10864 Segment
X10864 N10864 N10865 Segment
X10865 N10865 N10866 Segment
X10866 N10866 N10867 Segment
X10867 N10867 N10868 Segment
X10868 N10868 N10869 Segment
X10869 N10869 N10870 Segment
X10870 N10870 N10871 Segment
X10871 N10871 N10872 Segment
X10872 N10872 N10873 Segment
X10873 N10873 N10874 Segment
X10874 N10874 N10875 Segment
X10875 N10875 N10876 Segment
X10876 N10876 N10877 Segment
X10877 N10877 N10878 Segment
X10878 N10878 N10879 Segment
X10879 N10879 N10880 Segment
X10880 N10880 N10881 Segment
X10881 N10881 N10882 Segment
X10882 N10882 N10883 Segment
X10883 N10883 N10884 Segment
X10884 N10884 N10885 Segment
X10885 N10885 N10886 Segment
X10886 N10886 N10887 Segment
X10887 N10887 N10888 Segment
X10888 N10888 N10889 Segment
X10889 N10889 N10890 Segment
X10890 N10890 N10891 Segment
X10891 N10891 N10892 Segment
X10892 N10892 N10893 Segment
X10893 N10893 N10894 Segment
X10894 N10894 N10895 Segment
X10895 N10895 N10896 Segment
X10896 N10896 N10897 Segment
X10897 N10897 N10898 Segment
X10898 N10898 N10899 Segment
X10899 N10899 N10900 Segment
X10900 N10900 N10901 Segment
X10901 N10901 N10902 Segment
X10902 N10902 N10903 Segment
X10903 N10903 N10904 Segment
X10904 N10904 N10905 Segment
X10905 N10905 N10906 Segment
X10906 N10906 N10907 Segment
X10907 N10907 N10908 Segment
X10908 N10908 N10909 Segment
X10909 N10909 N10910 Segment
X10910 N10910 N10911 Segment
X10911 N10911 N10912 Segment
X10912 N10912 N10913 Segment
X10913 N10913 N10914 Segment
X10914 N10914 N10915 Segment
X10915 N10915 N10916 Segment
X10916 N10916 N10917 Segment
X10917 N10917 N10918 Segment
X10918 N10918 N10919 Segment
X10919 N10919 N10920 Segment
X10920 N10920 N10921 Segment
X10921 N10921 N10922 Segment
X10922 N10922 N10923 Segment
X10923 N10923 N10924 Segment
X10924 N10924 N10925 Segment
X10925 N10925 N10926 Segment
X10926 N10926 N10927 Segment
X10927 N10927 N10928 Segment
X10928 N10928 N10929 Segment
X10929 N10929 N10930 Segment
X10930 N10930 N10931 Segment
X10931 N10931 N10932 Segment
X10932 N10932 N10933 Segment
X10933 N10933 N10934 Segment
X10934 N10934 N10935 Segment
X10935 N10935 N10936 Segment
X10936 N10936 N10937 Segment
X10937 N10937 N10938 Segment
X10938 N10938 N10939 Segment
X10939 N10939 N10940 Segment
X10940 N10940 N10941 Segment
X10941 N10941 N10942 Segment
X10942 N10942 N10943 Segment
X10943 N10943 N10944 Segment
X10944 N10944 N10945 Segment
X10945 N10945 N10946 Segment
X10946 N10946 N10947 Segment
X10947 N10947 N10948 Segment
X10948 N10948 N10949 Segment
X10949 N10949 N10950 Segment
X10950 N10950 N10951 Segment
X10951 N10951 N10952 Segment
X10952 N10952 N10953 Segment
X10953 N10953 N10954 Segment
X10954 N10954 N10955 Segment
X10955 N10955 N10956 Segment
X10956 N10956 N10957 Segment
X10957 N10957 N10958 Segment
X10958 N10958 N10959 Segment
X10959 N10959 N10960 Segment
X10960 N10960 N10961 Segment
X10961 N10961 N10962 Segment
X10962 N10962 N10963 Segment
X10963 N10963 N10964 Segment
X10964 N10964 N10965 Segment
X10965 N10965 N10966 Segment
X10966 N10966 N10967 Segment
X10967 N10967 N10968 Segment
X10968 N10968 N10969 Segment
X10969 N10969 N10970 Segment
X10970 N10970 N10971 Segment
X10971 N10971 N10972 Segment
X10972 N10972 N10973 Segment
X10973 N10973 N10974 Segment
X10974 N10974 N10975 Segment
X10975 N10975 N10976 Segment
X10976 N10976 N10977 Segment
X10977 N10977 N10978 Segment
X10978 N10978 N10979 Segment
X10979 N10979 N10980 Segment
X10980 N10980 N10981 Segment
X10981 N10981 N10982 Segment
X10982 N10982 N10983 Segment
X10983 N10983 N10984 Segment
X10984 N10984 N10985 Segment
X10985 N10985 N10986 Segment
X10986 N10986 N10987 Segment
X10987 N10987 N10988 Segment
X10988 N10988 N10989 Segment
X10989 N10989 N10990 Segment
X10990 N10990 N10991 Segment
X10991 N10991 N10992 Segment
X10992 N10992 N10993 Segment
X10993 N10993 N10994 Segment
X10994 N10994 N10995 Segment
X10995 N10995 N10996 Segment
X10996 N10996 N10997 Segment
X10997 N10997 N10998 Segment
X10998 N10998 N10999 Segment
X10999 N10999 N11000 Segment
X11000 N11000 N11001 Segment
X11001 N11001 N11002 Segment
X11002 N11002 N11003 Segment
X11003 N11003 N11004 Segment
X11004 N11004 N11005 Segment
X11005 N11005 N11006 Segment
X11006 N11006 N11007 Segment
X11007 N11007 N11008 Segment
X11008 N11008 N11009 Segment
X11009 N11009 N11010 Segment
X11010 N11010 N11011 Segment
X11011 N11011 N11012 Segment
X11012 N11012 N11013 Segment
X11013 N11013 N11014 Segment
X11014 N11014 N11015 Segment
X11015 N11015 N11016 Segment
X11016 N11016 N11017 Segment
X11017 N11017 N11018 Segment
X11018 N11018 N11019 Segment
X11019 N11019 N11020 Segment
X11020 N11020 N11021 Segment
X11021 N11021 N11022 Segment
X11022 N11022 N11023 Segment
X11023 N11023 N11024 Segment
X11024 N11024 N11025 Segment
X11025 N11025 N11026 Segment
X11026 N11026 N11027 Segment
X11027 N11027 N11028 Segment
X11028 N11028 N11029 Segment
X11029 N11029 N11030 Segment
X11030 N11030 N11031 Segment
X11031 N11031 N11032 Segment
X11032 N11032 N11033 Segment
X11033 N11033 N11034 Segment
X11034 N11034 N11035 Segment
X11035 N11035 N11036 Segment
X11036 N11036 N11037 Segment
X11037 N11037 N11038 Segment
X11038 N11038 N11039 Segment
X11039 N11039 N11040 Segment
X11040 N11040 N11041 Segment
X11041 N11041 N11042 Segment
X11042 N11042 N11043 Segment
X11043 N11043 N11044 Segment
X11044 N11044 N11045 Segment
X11045 N11045 N11046 Segment
X11046 N11046 N11047 Segment
X11047 N11047 N11048 Segment
X11048 N11048 N11049 Segment
X11049 N11049 N11050 Segment
X11050 N11050 N11051 Segment
X11051 N11051 N11052 Segment
X11052 N11052 N11053 Segment
X11053 N11053 N11054 Segment
X11054 N11054 N11055 Segment
X11055 N11055 N11056 Segment
X11056 N11056 N11057 Segment
X11057 N11057 N11058 Segment
X11058 N11058 N11059 Segment
X11059 N11059 N11060 Segment
X11060 N11060 N11061 Segment
X11061 N11061 N11062 Segment
X11062 N11062 N11063 Segment
X11063 N11063 N11064 Segment
X11064 N11064 N11065 Segment
X11065 N11065 N11066 Segment
X11066 N11066 N11067 Segment
X11067 N11067 N11068 Segment
X11068 N11068 N11069 Segment
X11069 N11069 N11070 Segment
X11070 N11070 N11071 Segment
X11071 N11071 N11072 Segment
X11072 N11072 N11073 Segment
X11073 N11073 N11074 Segment
X11074 N11074 N11075 Segment
X11075 N11075 N11076 Segment
X11076 N11076 N11077 Segment
X11077 N11077 N11078 Segment
X11078 N11078 N11079 Segment
X11079 N11079 N11080 Segment
X11080 N11080 N11081 Segment
X11081 N11081 N11082 Segment
X11082 N11082 N11083 Segment
X11083 N11083 N11084 Segment
X11084 N11084 N11085 Segment
X11085 N11085 N11086 Segment
X11086 N11086 N11087 Segment
X11087 N11087 N11088 Segment
X11088 N11088 N11089 Segment
X11089 N11089 N11090 Segment
X11090 N11090 N11091 Segment
X11091 N11091 N11092 Segment
X11092 N11092 N11093 Segment
X11093 N11093 N11094 Segment
X11094 N11094 N11095 Segment
X11095 N11095 N11096 Segment
X11096 N11096 N11097 Segment
X11097 N11097 N11098 Segment
X11098 N11098 N11099 Segment
X11099 N11099 N11100 Segment
X11100 N11100 N11101 Segment
X11101 N11101 N11102 Segment
X11102 N11102 N11103 Segment
X11103 N11103 N11104 Segment
X11104 N11104 N11105 Segment
X11105 N11105 N11106 Segment
X11106 N11106 N11107 Segment
X11107 N11107 N11108 Segment
X11108 N11108 N11109 Segment
X11109 N11109 N11110 Segment
X11110 N11110 N11111 Segment
X11111 N11111 N11112 Segment
X11112 N11112 N11113 Segment
X11113 N11113 N11114 Segment
X11114 N11114 N11115 Segment
X11115 N11115 N11116 Segment
X11116 N11116 N11117 Segment
X11117 N11117 N11118 Segment
X11118 N11118 N11119 Segment
X11119 N11119 N11120 Segment
X11120 N11120 N11121 Segment
X11121 N11121 N11122 Segment
X11122 N11122 N11123 Segment
X11123 N11123 N11124 Segment
X11124 N11124 N11125 Segment
X11125 N11125 N11126 Segment
X11126 N11126 N11127 Segment
X11127 N11127 N11128 Segment
X11128 N11128 N11129 Segment
X11129 N11129 N11130 Segment
X11130 N11130 N11131 Segment
X11131 N11131 N11132 Segment
X11132 N11132 N11133 Segment
X11133 N11133 N11134 Segment
X11134 N11134 N11135 Segment
X11135 N11135 N11136 Segment
X11136 N11136 N11137 Segment
X11137 N11137 N11138 Segment
X11138 N11138 N11139 Segment
X11139 N11139 N11140 Segment
X11140 N11140 N11141 Segment
X11141 N11141 N11142 Segment
X11142 N11142 N11143 Segment
X11143 N11143 N11144 Segment
X11144 N11144 N11145 Segment
X11145 N11145 N11146 Segment
X11146 N11146 N11147 Segment
X11147 N11147 N11148 Segment
X11148 N11148 N11149 Segment
X11149 N11149 N11150 Segment
X11150 N11150 N11151 Segment
X11151 N11151 N11152 Segment
X11152 N11152 N11153 Segment
X11153 N11153 N11154 Segment
X11154 N11154 N11155 Segment
X11155 N11155 N11156 Segment
X11156 N11156 N11157 Segment
X11157 N11157 N11158 Segment
X11158 N11158 N11159 Segment
X11159 N11159 N11160 Segment
X11160 N11160 N11161 Segment
X11161 N11161 N11162 Segment
X11162 N11162 N11163 Segment
X11163 N11163 N11164 Segment
X11164 N11164 N11165 Segment
X11165 N11165 N11166 Segment
X11166 N11166 N11167 Segment
X11167 N11167 N11168 Segment
X11168 N11168 N11169 Segment
X11169 N11169 N11170 Segment
X11170 N11170 N11171 Segment
X11171 N11171 N11172 Segment
X11172 N11172 N11173 Segment
X11173 N11173 N11174 Segment
X11174 N11174 N11175 Segment
X11175 N11175 N11176 Segment
X11176 N11176 N11177 Segment
X11177 N11177 N11178 Segment
X11178 N11178 N11179 Segment
X11179 N11179 N11180 Segment
X11180 N11180 N11181 Segment
X11181 N11181 N11182 Segment
X11182 N11182 N11183 Segment
X11183 N11183 N11184 Segment
X11184 N11184 N11185 Segment
X11185 N11185 N11186 Segment
X11186 N11186 N11187 Segment
X11187 N11187 N11188 Segment
X11188 N11188 N11189 Segment
X11189 N11189 N11190 Segment
X11190 N11190 N11191 Segment
X11191 N11191 N11192 Segment
X11192 N11192 N11193 Segment
X11193 N11193 N11194 Segment
X11194 N11194 N11195 Segment
X11195 N11195 N11196 Segment
X11196 N11196 N11197 Segment
X11197 N11197 N11198 Segment
X11198 N11198 N11199 Segment
X11199 N11199 N11200 Segment
X11200 N11200 N11201 Segment
X11201 N11201 N11202 Segment
X11202 N11202 N11203 Segment
X11203 N11203 N11204 Segment
X11204 N11204 N11205 Segment
X11205 N11205 N11206 Segment
X11206 N11206 N11207 Segment
X11207 N11207 N11208 Segment
X11208 N11208 N11209 Segment
X11209 N11209 N11210 Segment
X11210 N11210 N11211 Segment
X11211 N11211 N11212 Segment
X11212 N11212 N11213 Segment
X11213 N11213 N11214 Segment
X11214 N11214 N11215 Segment
X11215 N11215 N11216 Segment
X11216 N11216 N11217 Segment
X11217 N11217 N11218 Segment
X11218 N11218 N11219 Segment
X11219 N11219 N11220 Segment
X11220 N11220 N11221 Segment
X11221 N11221 N11222 Segment
X11222 N11222 N11223 Segment
X11223 N11223 N11224 Segment
X11224 N11224 N11225 Segment
X11225 N11225 N11226 Segment
X11226 N11226 N11227 Segment
X11227 N11227 N11228 Segment
X11228 N11228 N11229 Segment
X11229 N11229 N11230 Segment
X11230 N11230 N11231 Segment
X11231 N11231 N11232 Segment
X11232 N11232 N11233 Segment
X11233 N11233 N11234 Segment
X11234 N11234 N11235 Segment
X11235 N11235 N11236 Segment
X11236 N11236 N11237 Segment
X11237 N11237 N11238 Segment
X11238 N11238 N11239 Segment
X11239 N11239 N11240 Segment
X11240 N11240 N11241 Segment
X11241 N11241 N11242 Segment
X11242 N11242 N11243 Segment
X11243 N11243 N11244 Segment
X11244 N11244 N11245 Segment
X11245 N11245 N11246 Segment
X11246 N11246 N11247 Segment
X11247 N11247 N11248 Segment
X11248 N11248 N11249 Segment
X11249 N11249 N11250 Segment
X11250 N11250 N11251 Segment
X11251 N11251 N11252 Segment
X11252 N11252 N11253 Segment
X11253 N11253 N11254 Segment
X11254 N11254 N11255 Segment
X11255 N11255 N11256 Segment
X11256 N11256 N11257 Segment
X11257 N11257 N11258 Segment
X11258 N11258 N11259 Segment
X11259 N11259 N11260 Segment
X11260 N11260 N11261 Segment
X11261 N11261 N11262 Segment
X11262 N11262 N11263 Segment
X11263 N11263 N11264 Segment
X11264 N11264 N11265 Segment
X11265 N11265 N11266 Segment
X11266 N11266 N11267 Segment
X11267 N11267 N11268 Segment
X11268 N11268 N11269 Segment
X11269 N11269 N11270 Segment
X11270 N11270 N11271 Segment
X11271 N11271 N11272 Segment
X11272 N11272 N11273 Segment
X11273 N11273 N11274 Segment
X11274 N11274 N11275 Segment
X11275 N11275 N11276 Segment
X11276 N11276 N11277 Segment
X11277 N11277 N11278 Segment
X11278 N11278 N11279 Segment
X11279 N11279 N11280 Segment
X11280 N11280 N11281 Segment
X11281 N11281 N11282 Segment
X11282 N11282 N11283 Segment
X11283 N11283 N11284 Segment
X11284 N11284 N11285 Segment
X11285 N11285 N11286 Segment
X11286 N11286 N11287 Segment
X11287 N11287 N11288 Segment
X11288 N11288 N11289 Segment
X11289 N11289 N11290 Segment
X11290 N11290 N11291 Segment
X11291 N11291 N11292 Segment
X11292 N11292 N11293 Segment
X11293 N11293 N11294 Segment
X11294 N11294 N11295 Segment
X11295 N11295 N11296 Segment
X11296 N11296 N11297 Segment
X11297 N11297 N11298 Segment
X11298 N11298 N11299 Segment
X11299 N11299 N11300 Segment
X11300 N11300 N11301 Segment
X11301 N11301 N11302 Segment
X11302 N11302 N11303 Segment
X11303 N11303 N11304 Segment
X11304 N11304 N11305 Segment
X11305 N11305 N11306 Segment
X11306 N11306 N11307 Segment
X11307 N11307 N11308 Segment
X11308 N11308 N11309 Segment
X11309 N11309 N11310 Segment
X11310 N11310 N11311 Segment
X11311 N11311 N11312 Segment
X11312 N11312 N11313 Segment
X11313 N11313 N11314 Segment
X11314 N11314 N11315 Segment
X11315 N11315 N11316 Segment
X11316 N11316 N11317 Segment
X11317 N11317 N11318 Segment
X11318 N11318 N11319 Segment
X11319 N11319 N11320 Segment
X11320 N11320 N11321 Segment
X11321 N11321 N11322 Segment
X11322 N11322 N11323 Segment
X11323 N11323 N11324 Segment
X11324 N11324 N11325 Segment
X11325 N11325 N11326 Segment
X11326 N11326 N11327 Segment
X11327 N11327 N11328 Segment
X11328 N11328 N11329 Segment
X11329 N11329 N11330 Segment
X11330 N11330 N11331 Segment
X11331 N11331 N11332 Segment
X11332 N11332 N11333 Segment
X11333 N11333 N11334 Segment
X11334 N11334 N11335 Segment
X11335 N11335 N11336 Segment
X11336 N11336 N11337 Segment
X11337 N11337 N11338 Segment
X11338 N11338 N11339 Segment
X11339 N11339 N11340 Segment
X11340 N11340 N11341 Segment
X11341 N11341 N11342 Segment
X11342 N11342 N11343 Segment
X11343 N11343 N11344 Segment
X11344 N11344 N11345 Segment
X11345 N11345 N11346 Segment
X11346 N11346 N11347 Segment
X11347 N11347 N11348 Segment
X11348 N11348 N11349 Segment
X11349 N11349 N11350 Segment
X11350 N11350 N11351 Segment
X11351 N11351 N11352 Segment
X11352 N11352 N11353 Segment
X11353 N11353 N11354 Segment
X11354 N11354 N11355 Segment
X11355 N11355 N11356 Segment
X11356 N11356 N11357 Segment
X11357 N11357 N11358 Segment
X11358 N11358 N11359 Segment
X11359 N11359 N11360 Segment
X11360 N11360 N11361 Segment
X11361 N11361 N11362 Segment
X11362 N11362 N11363 Segment
X11363 N11363 N11364 Segment
X11364 N11364 N11365 Segment
X11365 N11365 N11366 Segment
X11366 N11366 N11367 Segment
X11367 N11367 N11368 Segment
X11368 N11368 N11369 Segment
X11369 N11369 N11370 Segment
X11370 N11370 N11371 Segment
X11371 N11371 N11372 Segment
X11372 N11372 N11373 Segment
X11373 N11373 N11374 Segment
X11374 N11374 N11375 Segment
X11375 N11375 N11376 Segment
X11376 N11376 N11377 Segment
X11377 N11377 N11378 Segment
X11378 N11378 N11379 Segment
X11379 N11379 N11380 Segment
X11380 N11380 N11381 Segment
X11381 N11381 N11382 Segment
X11382 N11382 N11383 Segment
X11383 N11383 N11384 Segment
X11384 N11384 N11385 Segment
X11385 N11385 N11386 Segment
X11386 N11386 N11387 Segment
X11387 N11387 N11388 Segment
X11388 N11388 N11389 Segment
X11389 N11389 N11390 Segment
X11390 N11390 N11391 Segment
X11391 N11391 N11392 Segment
X11392 N11392 N11393 Segment
X11393 N11393 N11394 Segment
X11394 N11394 N11395 Segment
X11395 N11395 N11396 Segment
X11396 N11396 N11397 Segment
X11397 N11397 N11398 Segment
X11398 N11398 N11399 Segment
X11399 N11399 N11400 Segment
X11400 N11400 N11401 Segment
X11401 N11401 N11402 Segment
X11402 N11402 N11403 Segment
X11403 N11403 N11404 Segment
X11404 N11404 N11405 Segment
X11405 N11405 N11406 Segment
X11406 N11406 N11407 Segment
X11407 N11407 N11408 Segment
X11408 N11408 N11409 Segment
X11409 N11409 N11410 Segment
X11410 N11410 N11411 Segment
X11411 N11411 N11412 Segment
X11412 N11412 N11413 Segment
X11413 N11413 N11414 Segment
X11414 N11414 N11415 Segment
X11415 N11415 N11416 Segment
X11416 N11416 N11417 Segment
X11417 N11417 N11418 Segment
X11418 N11418 N11419 Segment
X11419 N11419 N11420 Segment
X11420 N11420 N11421 Segment
X11421 N11421 N11422 Segment
X11422 N11422 N11423 Segment
X11423 N11423 N11424 Segment
X11424 N11424 N11425 Segment
X11425 N11425 N11426 Segment
X11426 N11426 N11427 Segment
X11427 N11427 N11428 Segment
X11428 N11428 N11429 Segment
X11429 N11429 N11430 Segment
X11430 N11430 N11431 Segment
X11431 N11431 N11432 Segment
X11432 N11432 N11433 Segment
X11433 N11433 N11434 Segment
X11434 N11434 N11435 Segment
X11435 N11435 N11436 Segment
X11436 N11436 N11437 Segment
X11437 N11437 N11438 Segment
X11438 N11438 N11439 Segment
X11439 N11439 N11440 Segment
X11440 N11440 N11441 Segment
X11441 N11441 N11442 Segment
X11442 N11442 N11443 Segment
X11443 N11443 N11444 Segment
X11444 N11444 N11445 Segment
X11445 N11445 N11446 Segment
X11446 N11446 N11447 Segment
X11447 N11447 N11448 Segment
X11448 N11448 N11449 Segment
X11449 N11449 N11450 Segment
X11450 N11450 N11451 Segment
X11451 N11451 N11452 Segment
X11452 N11452 N11453 Segment
X11453 N11453 N11454 Segment
X11454 N11454 N11455 Segment
X11455 N11455 N11456 Segment
X11456 N11456 N11457 Segment
X11457 N11457 N11458 Segment
X11458 N11458 N11459 Segment
X11459 N11459 N11460 Segment
X11460 N11460 N11461 Segment
X11461 N11461 N11462 Segment
X11462 N11462 N11463 Segment
X11463 N11463 N11464 Segment
X11464 N11464 N11465 Segment
X11465 N11465 N11466 Segment
X11466 N11466 N11467 Segment
X11467 N11467 N11468 Segment
X11468 N11468 N11469 Segment
X11469 N11469 N11470 Segment
X11470 N11470 N11471 Segment
X11471 N11471 N11472 Segment
X11472 N11472 N11473 Segment
X11473 N11473 N11474 Segment
X11474 N11474 N11475 Segment
X11475 N11475 N11476 Segment
X11476 N11476 N11477 Segment
X11477 N11477 N11478 Segment
X11478 N11478 N11479 Segment
X11479 N11479 N11480 Segment
X11480 N11480 N11481 Segment
X11481 N11481 N11482 Segment
X11482 N11482 N11483 Segment
X11483 N11483 N11484 Segment
X11484 N11484 N11485 Segment
X11485 N11485 N11486 Segment
X11486 N11486 N11487 Segment
X11487 N11487 N11488 Segment
X11488 N11488 N11489 Segment
X11489 N11489 N11490 Segment
X11490 N11490 N11491 Segment
X11491 N11491 N11492 Segment
X11492 N11492 N11493 Segment
X11493 N11493 N11494 Segment
X11494 N11494 N11495 Segment
X11495 N11495 N11496 Segment
X11496 N11496 N11497 Segment
X11497 N11497 N11498 Segment
X11498 N11498 N11499 Segment
X11499 N11499 N11500 Segment
X11500 N11500 N11501 Segment
X11501 N11501 N11502 Segment
X11502 N11502 N11503 Segment
X11503 N11503 N11504 Segment
X11504 N11504 N11505 Segment
X11505 N11505 N11506 Segment
X11506 N11506 N11507 Segment
X11507 N11507 N11508 Segment
X11508 N11508 N11509 Segment
X11509 N11509 N11510 Segment
X11510 N11510 N11511 Segment
X11511 N11511 N11512 Segment
X11512 N11512 N11513 Segment
X11513 N11513 N11514 Segment
X11514 N11514 N11515 Segment
X11515 N11515 N11516 Segment
X11516 N11516 N11517 Segment
X11517 N11517 N11518 Segment
X11518 N11518 N11519 Segment
X11519 N11519 N11520 Segment
X11520 N11520 N11521 Segment
X11521 N11521 N11522 Segment
X11522 N11522 N11523 Segment
X11523 N11523 N11524 Segment
X11524 N11524 N11525 Segment
X11525 N11525 N11526 Segment
X11526 N11526 N11527 Segment
X11527 N11527 N11528 Segment
X11528 N11528 N11529 Segment
X11529 N11529 N11530 Segment
X11530 N11530 N11531 Segment
X11531 N11531 N11532 Segment
X11532 N11532 N11533 Segment
X11533 N11533 N11534 Segment
X11534 N11534 N11535 Segment
X11535 N11535 N11536 Segment
X11536 N11536 N11537 Segment
X11537 N11537 N11538 Segment
X11538 N11538 N11539 Segment
X11539 N11539 N11540 Segment
X11540 N11540 N11541 Segment
X11541 N11541 N11542 Segment
X11542 N11542 N11543 Segment
X11543 N11543 N11544 Segment
X11544 N11544 N11545 Segment
X11545 N11545 N11546 Segment
X11546 N11546 N11547 Segment
X11547 N11547 N11548 Segment
X11548 N11548 N11549 Segment
X11549 N11549 N11550 Segment
X11550 N11550 N11551 Segment
X11551 N11551 N11552 Segment
X11552 N11552 N11553 Segment
X11553 N11553 N11554 Segment
X11554 N11554 N11555 Segment
X11555 N11555 N11556 Segment
X11556 N11556 N11557 Segment
X11557 N11557 N11558 Segment
X11558 N11558 N11559 Segment
X11559 N11559 N11560 Segment
X11560 N11560 N11561 Segment
X11561 N11561 N11562 Segment
X11562 N11562 N11563 Segment
X11563 N11563 N11564 Segment
X11564 N11564 N11565 Segment
X11565 N11565 N11566 Segment
X11566 N11566 N11567 Segment
X11567 N11567 N11568 Segment
X11568 N11568 N11569 Segment
X11569 N11569 N11570 Segment
X11570 N11570 N11571 Segment
X11571 N11571 N11572 Segment
X11572 N11572 N11573 Segment
X11573 N11573 N11574 Segment
X11574 N11574 N11575 Segment
X11575 N11575 N11576 Segment
X11576 N11576 N11577 Segment
X11577 N11577 N11578 Segment
X11578 N11578 N11579 Segment
X11579 N11579 N11580 Segment
X11580 N11580 N11581 Segment
X11581 N11581 N11582 Segment
X11582 N11582 N11583 Segment
X11583 N11583 N11584 Segment
X11584 N11584 N11585 Segment
X11585 N11585 N11586 Segment
X11586 N11586 N11587 Segment
X11587 N11587 N11588 Segment
X11588 N11588 N11589 Segment
X11589 N11589 N11590 Segment
X11590 N11590 N11591 Segment
X11591 N11591 N11592 Segment
X11592 N11592 N11593 Segment
X11593 N11593 N11594 Segment
X11594 N11594 N11595 Segment
X11595 N11595 N11596 Segment
X11596 N11596 N11597 Segment
X11597 N11597 N11598 Segment
X11598 N11598 N11599 Segment
X11599 N11599 N11600 Segment
X11600 N11600 N11601 Segment
X11601 N11601 N11602 Segment
X11602 N11602 N11603 Segment
X11603 N11603 N11604 Segment
X11604 N11604 N11605 Segment
X11605 N11605 N11606 Segment
X11606 N11606 N11607 Segment
X11607 N11607 N11608 Segment
X11608 N11608 N11609 Segment
X11609 N11609 N11610 Segment
X11610 N11610 N11611 Segment
X11611 N11611 N11612 Segment
X11612 N11612 N11613 Segment
X11613 N11613 N11614 Segment
X11614 N11614 N11615 Segment
X11615 N11615 N11616 Segment
X11616 N11616 N11617 Segment
X11617 N11617 N11618 Segment
X11618 N11618 N11619 Segment
X11619 N11619 N11620 Segment
X11620 N11620 N11621 Segment
X11621 N11621 N11622 Segment
X11622 N11622 N11623 Segment
X11623 N11623 N11624 Segment
X11624 N11624 N11625 Segment
X11625 N11625 N11626 Segment
X11626 N11626 N11627 Segment
X11627 N11627 N11628 Segment
X11628 N11628 N11629 Segment
X11629 N11629 N11630 Segment
X11630 N11630 N11631 Segment
X11631 N11631 N11632 Segment
X11632 N11632 N11633 Segment
X11633 N11633 N11634 Segment
X11634 N11634 N11635 Segment
X11635 N11635 N11636 Segment
X11636 N11636 N11637 Segment
X11637 N11637 N11638 Segment
X11638 N11638 N11639 Segment
X11639 N11639 N11640 Segment
X11640 N11640 N11641 Segment
X11641 N11641 N11642 Segment
X11642 N11642 N11643 Segment
X11643 N11643 N11644 Segment
X11644 N11644 N11645 Segment
X11645 N11645 N11646 Segment
X11646 N11646 N11647 Segment
X11647 N11647 N11648 Segment
X11648 N11648 N11649 Segment
X11649 N11649 N11650 Segment
X11650 N11650 N11651 Segment
X11651 N11651 N11652 Segment
X11652 N11652 N11653 Segment
X11653 N11653 N11654 Segment
X11654 N11654 N11655 Segment
X11655 N11655 N11656 Segment
X11656 N11656 N11657 Segment
X11657 N11657 N11658 Segment
X11658 N11658 N11659 Segment
X11659 N11659 N11660 Segment
X11660 N11660 N11661 Segment
X11661 N11661 N11662 Segment
X11662 N11662 N11663 Segment
X11663 N11663 N11664 Segment
X11664 N11664 N11665 Segment
X11665 N11665 N11666 Segment
X11666 N11666 N11667 Segment
X11667 N11667 N11668 Segment
X11668 N11668 N11669 Segment
X11669 N11669 N11670 Segment
X11670 N11670 N11671 Segment
X11671 N11671 N11672 Segment
X11672 N11672 N11673 Segment
X11673 N11673 N11674 Segment
X11674 N11674 N11675 Segment
X11675 N11675 N11676 Segment
X11676 N11676 N11677 Segment
X11677 N11677 N11678 Segment
X11678 N11678 N11679 Segment
X11679 N11679 N11680 Segment
X11680 N11680 N11681 Segment
X11681 N11681 N11682 Segment
X11682 N11682 N11683 Segment
X11683 N11683 N11684 Segment
X11684 N11684 N11685 Segment
X11685 N11685 N11686 Segment
X11686 N11686 N11687 Segment
X11687 N11687 N11688 Segment
X11688 N11688 N11689 Segment
X11689 N11689 N11690 Segment
X11690 N11690 N11691 Segment
X11691 N11691 N11692 Segment
X11692 N11692 N11693 Segment
X11693 N11693 N11694 Segment
X11694 N11694 N11695 Segment
X11695 N11695 N11696 Segment
X11696 N11696 N11697 Segment
X11697 N11697 N11698 Segment
X11698 N11698 N11699 Segment
X11699 N11699 N11700 Segment
X11700 N11700 N11701 Segment
X11701 N11701 N11702 Segment
X11702 N11702 N11703 Segment
X11703 N11703 N11704 Segment
X11704 N11704 N11705 Segment
X11705 N11705 N11706 Segment
X11706 N11706 N11707 Segment
X11707 N11707 N11708 Segment
X11708 N11708 N11709 Segment
X11709 N11709 N11710 Segment
X11710 N11710 N11711 Segment
X11711 N11711 N11712 Segment
X11712 N11712 N11713 Segment
X11713 N11713 N11714 Segment
X11714 N11714 N11715 Segment
X11715 N11715 N11716 Segment
X11716 N11716 N11717 Segment
X11717 N11717 N11718 Segment
X11718 N11718 N11719 Segment
X11719 N11719 N11720 Segment
X11720 N11720 N11721 Segment
X11721 N11721 N11722 Segment
X11722 N11722 N11723 Segment
X11723 N11723 N11724 Segment
X11724 N11724 N11725 Segment
X11725 N11725 N11726 Segment
X11726 N11726 N11727 Segment
X11727 N11727 N11728 Segment
X11728 N11728 N11729 Segment
X11729 N11729 N11730 Segment
X11730 N11730 N11731 Segment
X11731 N11731 N11732 Segment
X11732 N11732 N11733 Segment
X11733 N11733 N11734 Segment
X11734 N11734 N11735 Segment
X11735 N11735 N11736 Segment
X11736 N11736 N11737 Segment
X11737 N11737 N11738 Segment
X11738 N11738 N11739 Segment
X11739 N11739 N11740 Segment
X11740 N11740 N11741 Segment
X11741 N11741 N11742 Segment
X11742 N11742 N11743 Segment
X11743 N11743 N11744 Segment
X11744 N11744 N11745 Segment
X11745 N11745 N11746 Segment
X11746 N11746 N11747 Segment
X11747 N11747 N11748 Segment
X11748 N11748 N11749 Segment
X11749 N11749 N11750 Segment
X11750 N11750 N11751 Segment
X11751 N11751 N11752 Segment
X11752 N11752 N11753 Segment
X11753 N11753 N11754 Segment
X11754 N11754 N11755 Segment
X11755 N11755 N11756 Segment
X11756 N11756 N11757 Segment
X11757 N11757 N11758 Segment
X11758 N11758 N11759 Segment
X11759 N11759 N11760 Segment
X11760 N11760 N11761 Segment
X11761 N11761 N11762 Segment
X11762 N11762 N11763 Segment
X11763 N11763 N11764 Segment
X11764 N11764 N11765 Segment
X11765 N11765 N11766 Segment
X11766 N11766 N11767 Segment
X11767 N11767 N11768 Segment
X11768 N11768 N11769 Segment
X11769 N11769 N11770 Segment
X11770 N11770 N11771 Segment
X11771 N11771 N11772 Segment
X11772 N11772 N11773 Segment
X11773 N11773 N11774 Segment
X11774 N11774 N11775 Segment
X11775 N11775 N11776 Segment
X11776 N11776 N11777 Segment
X11777 N11777 N11778 Segment
X11778 N11778 N11779 Segment
X11779 N11779 N11780 Segment
X11780 N11780 N11781 Segment
X11781 N11781 N11782 Segment
X11782 N11782 N11783 Segment
X11783 N11783 N11784 Segment
X11784 N11784 N11785 Segment
X11785 N11785 N11786 Segment
X11786 N11786 N11787 Segment
X11787 N11787 N11788 Segment
X11788 N11788 N11789 Segment
X11789 N11789 N11790 Segment
X11790 N11790 N11791 Segment
X11791 N11791 N11792 Segment
X11792 N11792 N11793 Segment
X11793 N11793 N11794 Segment
X11794 N11794 N11795 Segment
X11795 N11795 N11796 Segment
X11796 N11796 N11797 Segment
X11797 N11797 N11798 Segment
X11798 N11798 N11799 Segment
X11799 N11799 N11800 Segment
X11800 N11800 N11801 Segment
X11801 N11801 N11802 Segment
X11802 N11802 N11803 Segment
X11803 N11803 N11804 Segment
X11804 N11804 N11805 Segment
X11805 N11805 N11806 Segment
X11806 N11806 N11807 Segment
X11807 N11807 N11808 Segment
X11808 N11808 N11809 Segment
X11809 N11809 N11810 Segment
X11810 N11810 N11811 Segment
X11811 N11811 N11812 Segment
X11812 N11812 N11813 Segment
X11813 N11813 N11814 Segment
X11814 N11814 N11815 Segment
X11815 N11815 N11816 Segment
X11816 N11816 N11817 Segment
X11817 N11817 N11818 Segment
X11818 N11818 N11819 Segment
X11819 N11819 N11820 Segment
X11820 N11820 N11821 Segment
X11821 N11821 N11822 Segment
X11822 N11822 N11823 Segment
X11823 N11823 N11824 Segment
X11824 N11824 N11825 Segment
X11825 N11825 N11826 Segment
X11826 N11826 N11827 Segment
X11827 N11827 N11828 Segment
X11828 N11828 N11829 Segment
X11829 N11829 N11830 Segment
X11830 N11830 N11831 Segment
X11831 N11831 N11832 Segment
X11832 N11832 N11833 Segment
X11833 N11833 N11834 Segment
X11834 N11834 N11835 Segment
X11835 N11835 N11836 Segment
X11836 N11836 N11837 Segment
X11837 N11837 N11838 Segment
X11838 N11838 N11839 Segment
X11839 N11839 N11840 Segment
X11840 N11840 N11841 Segment
X11841 N11841 N11842 Segment
X11842 N11842 N11843 Segment
X11843 N11843 N11844 Segment
X11844 N11844 N11845 Segment
X11845 N11845 N11846 Segment
X11846 N11846 N11847 Segment
X11847 N11847 N11848 Segment
X11848 N11848 N11849 Segment
X11849 N11849 N11850 Segment
X11850 N11850 N11851 Segment
X11851 N11851 N11852 Segment
X11852 N11852 N11853 Segment
X11853 N11853 N11854 Segment
X11854 N11854 N11855 Segment
X11855 N11855 N11856 Segment
X11856 N11856 N11857 Segment
X11857 N11857 N11858 Segment
X11858 N11858 N11859 Segment
X11859 N11859 N11860 Segment
X11860 N11860 N11861 Segment
X11861 N11861 N11862 Segment
X11862 N11862 N11863 Segment
X11863 N11863 N11864 Segment
X11864 N11864 N11865 Segment
X11865 N11865 N11866 Segment
X11866 N11866 N11867 Segment
X11867 N11867 N11868 Segment
X11868 N11868 N11869 Segment
X11869 N11869 N11870 Segment
X11870 N11870 N11871 Segment
X11871 N11871 N11872 Segment
X11872 N11872 N11873 Segment
X11873 N11873 N11874 Segment
X11874 N11874 N11875 Segment
X11875 N11875 N11876 Segment
X11876 N11876 N11877 Segment
X11877 N11877 N11878 Segment
X11878 N11878 N11879 Segment
X11879 N11879 N11880 Segment
X11880 N11880 N11881 Segment
X11881 N11881 N11882 Segment
X11882 N11882 N11883 Segment
X11883 N11883 N11884 Segment
X11884 N11884 N11885 Segment
X11885 N11885 N11886 Segment
X11886 N11886 N11887 Segment
X11887 N11887 N11888 Segment
X11888 N11888 N11889 Segment
X11889 N11889 N11890 Segment
X11890 N11890 N11891 Segment
X11891 N11891 N11892 Segment
X11892 N11892 N11893 Segment
X11893 N11893 N11894 Segment
X11894 N11894 N11895 Segment
X11895 N11895 N11896 Segment
X11896 N11896 N11897 Segment
X11897 N11897 N11898 Segment
X11898 N11898 N11899 Segment
X11899 N11899 N11900 Segment
X11900 N11900 N11901 Segment
X11901 N11901 N11902 Segment
X11902 N11902 N11903 Segment
X11903 N11903 N11904 Segment
X11904 N11904 N11905 Segment
X11905 N11905 N11906 Segment
X11906 N11906 N11907 Segment
X11907 N11907 N11908 Segment
X11908 N11908 N11909 Segment
X11909 N11909 N11910 Segment
X11910 N11910 N11911 Segment
X11911 N11911 N11912 Segment
X11912 N11912 N11913 Segment
X11913 N11913 N11914 Segment
X11914 N11914 N11915 Segment
X11915 N11915 N11916 Segment
X11916 N11916 N11917 Segment
X11917 N11917 N11918 Segment
X11918 N11918 N11919 Segment
X11919 N11919 N11920 Segment
X11920 N11920 N11921 Segment
X11921 N11921 N11922 Segment
X11922 N11922 N11923 Segment
X11923 N11923 N11924 Segment
X11924 N11924 N11925 Segment
X11925 N11925 N11926 Segment
X11926 N11926 N11927 Segment
X11927 N11927 N11928 Segment
X11928 N11928 N11929 Segment
X11929 N11929 N11930 Segment
X11930 N11930 N11931 Segment
X11931 N11931 N11932 Segment
X11932 N11932 N11933 Segment
X11933 N11933 N11934 Segment
X11934 N11934 N11935 Segment
X11935 N11935 N11936 Segment
X11936 N11936 N11937 Segment
X11937 N11937 N11938 Segment
X11938 N11938 N11939 Segment
X11939 N11939 N11940 Segment
X11940 N11940 N11941 Segment
X11941 N11941 N11942 Segment
X11942 N11942 N11943 Segment
X11943 N11943 N11944 Segment
X11944 N11944 N11945 Segment
X11945 N11945 N11946 Segment
X11946 N11946 N11947 Segment
X11947 N11947 N11948 Segment
X11948 N11948 N11949 Segment
X11949 N11949 N11950 Segment
X11950 N11950 N11951 Segment
X11951 N11951 N11952 Segment
X11952 N11952 N11953 Segment
X11953 N11953 N11954 Segment
X11954 N11954 N11955 Segment
X11955 N11955 N11956 Segment
X11956 N11956 N11957 Segment
X11957 N11957 N11958 Segment
X11958 N11958 N11959 Segment
X11959 N11959 N11960 Segment
X11960 N11960 N11961 Segment
X11961 N11961 N11962 Segment
X11962 N11962 N11963 Segment
X11963 N11963 N11964 Segment
X11964 N11964 N11965 Segment
X11965 N11965 N11966 Segment
X11966 N11966 N11967 Segment
X11967 N11967 N11968 Segment
X11968 N11968 N11969 Segment
X11969 N11969 N11970 Segment
X11970 N11970 N11971 Segment
X11971 N11971 N11972 Segment
X11972 N11972 N11973 Segment
X11973 N11973 N11974 Segment
X11974 N11974 N11975 Segment
X11975 N11975 N11976 Segment
X11976 N11976 N11977 Segment
X11977 N11977 N11978 Segment
X11978 N11978 N11979 Segment
X11979 N11979 N11980 Segment
X11980 N11980 N11981 Segment
X11981 N11981 N11982 Segment
X11982 N11982 N11983 Segment
X11983 N11983 N11984 Segment
X11984 N11984 N11985 Segment
X11985 N11985 N11986 Segment
X11986 N11986 N11987 Segment
X11987 N11987 N11988 Segment
X11988 N11988 N11989 Segment
X11989 N11989 N11990 Segment
X11990 N11990 N11991 Segment
X11991 N11991 N11992 Segment
X11992 N11992 N11993 Segment
X11993 N11993 N11994 Segment
X11994 N11994 N11995 Segment
X11995 N11995 N11996 Segment
X11996 N11996 N11997 Segment
X11997 N11997 N11998 Segment
X11998 N11998 N11999 Segment
X11999 N11999 N12000 Segment
X12000 N12000 N12001 Segment
X12001 N12001 N12002 Segment
X12002 N12002 N12003 Segment
X12003 N12003 N12004 Segment
X12004 N12004 N12005 Segment
X12005 N12005 N12006 Segment
X12006 N12006 N12007 Segment
X12007 N12007 N12008 Segment
X12008 N12008 N12009 Segment
X12009 N12009 N12010 Segment
X12010 N12010 N12011 Segment
X12011 N12011 N12012 Segment
X12012 N12012 N12013 Segment
X12013 N12013 N12014 Segment
X12014 N12014 N12015 Segment
X12015 N12015 N12016 Segment
X12016 N12016 N12017 Segment
X12017 N12017 N12018 Segment
X12018 N12018 N12019 Segment
X12019 N12019 N12020 Segment
X12020 N12020 N12021 Segment
X12021 N12021 N12022 Segment
X12022 N12022 N12023 Segment
X12023 N12023 N12024 Segment
X12024 N12024 N12025 Segment
X12025 N12025 N12026 Segment
X12026 N12026 N12027 Segment
X12027 N12027 N12028 Segment
X12028 N12028 N12029 Segment
X12029 N12029 N12030 Segment
X12030 N12030 N12031 Segment
X12031 N12031 N12032 Segment
X12032 N12032 N12033 Segment
X12033 N12033 N12034 Segment
X12034 N12034 N12035 Segment
X12035 N12035 N12036 Segment
X12036 N12036 N12037 Segment
X12037 N12037 N12038 Segment
X12038 N12038 N12039 Segment
X12039 N12039 N12040 Segment
X12040 N12040 N12041 Segment
X12041 N12041 N12042 Segment
X12042 N12042 N12043 Segment
X12043 N12043 N12044 Segment
X12044 N12044 N12045 Segment
X12045 N12045 N12046 Segment
X12046 N12046 N12047 Segment
X12047 N12047 N12048 Segment
X12048 N12048 N12049 Segment
X12049 N12049 N12050 Segment
X12050 N12050 N12051 Segment
X12051 N12051 N12052 Segment
X12052 N12052 N12053 Segment
X12053 N12053 N12054 Segment
X12054 N12054 N12055 Segment
X12055 N12055 N12056 Segment
X12056 N12056 N12057 Segment
X12057 N12057 N12058 Segment
X12058 N12058 N12059 Segment
X12059 N12059 N12060 Segment
X12060 N12060 N12061 Segment
X12061 N12061 N12062 Segment
X12062 N12062 N12063 Segment
X12063 N12063 N12064 Segment
X12064 N12064 N12065 Segment
X12065 N12065 N12066 Segment
X12066 N12066 N12067 Segment
X12067 N12067 N12068 Segment
X12068 N12068 N12069 Segment
X12069 N12069 N12070 Segment
X12070 N12070 N12071 Segment
X12071 N12071 N12072 Segment
X12072 N12072 N12073 Segment
X12073 N12073 N12074 Segment
X12074 N12074 N12075 Segment
X12075 N12075 N12076 Segment
X12076 N12076 N12077 Segment
X12077 N12077 N12078 Segment
X12078 N12078 N12079 Segment
X12079 N12079 N12080 Segment
X12080 N12080 N12081 Segment
X12081 N12081 N12082 Segment
X12082 N12082 N12083 Segment
X12083 N12083 N12084 Segment
X12084 N12084 N12085 Segment
X12085 N12085 N12086 Segment
X12086 N12086 N12087 Segment
X12087 N12087 N12088 Segment
X12088 N12088 N12089 Segment
X12089 N12089 N12090 Segment
X12090 N12090 N12091 Segment
X12091 N12091 N12092 Segment
X12092 N12092 N12093 Segment
X12093 N12093 N12094 Segment
X12094 N12094 N12095 Segment
X12095 N12095 N12096 Segment
X12096 N12096 N12097 Segment
X12097 N12097 N12098 Segment
X12098 N12098 N12099 Segment
X12099 N12099 N12100 Segment
X12100 N12100 N12101 Segment
X12101 N12101 N12102 Segment
X12102 N12102 N12103 Segment
X12103 N12103 N12104 Segment
X12104 N12104 N12105 Segment
X12105 N12105 N12106 Segment
X12106 N12106 N12107 Segment
X12107 N12107 N12108 Segment
X12108 N12108 N12109 Segment
X12109 N12109 N12110 Segment
X12110 N12110 N12111 Segment
X12111 N12111 N12112 Segment
X12112 N12112 N12113 Segment
X12113 N12113 N12114 Segment
X12114 N12114 N12115 Segment
X12115 N12115 N12116 Segment
X12116 N12116 N12117 Segment
X12117 N12117 N12118 Segment
X12118 N12118 N12119 Segment
X12119 N12119 N12120 Segment
X12120 N12120 N12121 Segment
X12121 N12121 N12122 Segment
X12122 N12122 N12123 Segment
X12123 N12123 N12124 Segment
X12124 N12124 N12125 Segment
X12125 N12125 N12126 Segment
X12126 N12126 N12127 Segment
X12127 N12127 N12128 Segment
X12128 N12128 N12129 Segment
X12129 N12129 N12130 Segment
X12130 N12130 N12131 Segment
X12131 N12131 N12132 Segment
X12132 N12132 N12133 Segment
X12133 N12133 N12134 Segment
X12134 N12134 N12135 Segment
X12135 N12135 N12136 Segment
X12136 N12136 N12137 Segment
X12137 N12137 N12138 Segment
X12138 N12138 N12139 Segment
X12139 N12139 N12140 Segment
X12140 N12140 N12141 Segment
X12141 N12141 N12142 Segment
X12142 N12142 N12143 Segment
X12143 N12143 N12144 Segment
X12144 N12144 N12145 Segment
X12145 N12145 N12146 Segment
X12146 N12146 N12147 Segment
X12147 N12147 N12148 Segment
X12148 N12148 N12149 Segment
X12149 N12149 N12150 Segment
X12150 N12150 N12151 Segment
X12151 N12151 N12152 Segment
X12152 N12152 N12153 Segment
X12153 N12153 N12154 Segment
X12154 N12154 N12155 Segment
X12155 N12155 N12156 Segment
X12156 N12156 N12157 Segment
X12157 N12157 N12158 Segment
X12158 N12158 N12159 Segment
X12159 N12159 N12160 Segment
X12160 N12160 N12161 Segment
X12161 N12161 N12162 Segment
X12162 N12162 N12163 Segment
X12163 N12163 N12164 Segment
X12164 N12164 N12165 Segment
X12165 N12165 N12166 Segment
X12166 N12166 N12167 Segment
X12167 N12167 N12168 Segment
X12168 N12168 N12169 Segment
X12169 N12169 N12170 Segment
X12170 N12170 N12171 Segment
X12171 N12171 N12172 Segment
X12172 N12172 N12173 Segment
X12173 N12173 N12174 Segment
X12174 N12174 N12175 Segment
X12175 N12175 N12176 Segment
X12176 N12176 N12177 Segment
X12177 N12177 N12178 Segment
X12178 N12178 N12179 Segment
X12179 N12179 N12180 Segment
X12180 N12180 N12181 Segment
X12181 N12181 N12182 Segment
X12182 N12182 N12183 Segment
X12183 N12183 N12184 Segment
X12184 N12184 N12185 Segment
X12185 N12185 N12186 Segment
X12186 N12186 N12187 Segment
X12187 N12187 N12188 Segment
X12188 N12188 N12189 Segment
X12189 N12189 N12190 Segment
X12190 N12190 N12191 Segment
X12191 N12191 N12192 Segment
X12192 N12192 N12193 Segment
X12193 N12193 N12194 Segment
X12194 N12194 N12195 Segment
X12195 N12195 N12196 Segment
X12196 N12196 N12197 Segment
X12197 N12197 N12198 Segment
X12198 N12198 N12199 Segment
X12199 N12199 N12200 Segment
X12200 N12200 N12201 Segment
X12201 N12201 N12202 Segment
X12202 N12202 N12203 Segment
X12203 N12203 N12204 Segment
X12204 N12204 N12205 Segment
X12205 N12205 N12206 Segment
X12206 N12206 N12207 Segment
X12207 N12207 N12208 Segment
X12208 N12208 N12209 Segment
X12209 N12209 N12210 Segment
X12210 N12210 N12211 Segment
X12211 N12211 N12212 Segment
X12212 N12212 N12213 Segment
X12213 N12213 N12214 Segment
X12214 N12214 N12215 Segment
X12215 N12215 N12216 Segment
X12216 N12216 N12217 Segment
X12217 N12217 N12218 Segment
X12218 N12218 N12219 Segment
X12219 N12219 N12220 Segment
X12220 N12220 N12221 Segment
X12221 N12221 N12222 Segment
X12222 N12222 N12223 Segment
X12223 N12223 N12224 Segment
X12224 N12224 N12225 Segment
X12225 N12225 N12226 Segment
X12226 N12226 N12227 Segment
X12227 N12227 N12228 Segment
X12228 N12228 N12229 Segment
X12229 N12229 N12230 Segment
X12230 N12230 N12231 Segment
X12231 N12231 N12232 Segment
X12232 N12232 N12233 Segment
X12233 N12233 N12234 Segment
X12234 N12234 N12235 Segment
X12235 N12235 N12236 Segment
X12236 N12236 N12237 Segment
X12237 N12237 N12238 Segment
X12238 N12238 N12239 Segment
X12239 N12239 N12240 Segment
X12240 N12240 N12241 Segment
X12241 N12241 N12242 Segment
X12242 N12242 N12243 Segment
X12243 N12243 N12244 Segment
X12244 N12244 N12245 Segment
X12245 N12245 N12246 Segment
X12246 N12246 N12247 Segment
X12247 N12247 N12248 Segment
X12248 N12248 N12249 Segment
X12249 N12249 N12250 Segment
X12250 N12250 N12251 Segment
X12251 N12251 N12252 Segment
X12252 N12252 N12253 Segment
X12253 N12253 N12254 Segment
X12254 N12254 N12255 Segment
X12255 N12255 N12256 Segment
X12256 N12256 N12257 Segment
X12257 N12257 N12258 Segment
X12258 N12258 N12259 Segment
X12259 N12259 N12260 Segment
X12260 N12260 N12261 Segment
X12261 N12261 N12262 Segment
X12262 N12262 N12263 Segment
X12263 N12263 N12264 Segment
X12264 N12264 N12265 Segment
X12265 N12265 N12266 Segment
X12266 N12266 N12267 Segment
X12267 N12267 N12268 Segment
X12268 N12268 N12269 Segment
X12269 N12269 N12270 Segment
X12270 N12270 N12271 Segment
X12271 N12271 N12272 Segment
X12272 N12272 N12273 Segment
X12273 N12273 N12274 Segment
X12274 N12274 N12275 Segment
X12275 N12275 N12276 Segment
X12276 N12276 N12277 Segment
X12277 N12277 N12278 Segment
X12278 N12278 N12279 Segment
X12279 N12279 N12280 Segment
X12280 N12280 N12281 Segment
X12281 N12281 N12282 Segment
X12282 N12282 N12283 Segment
X12283 N12283 N12284 Segment
X12284 N12284 N12285 Segment
X12285 N12285 N12286 Segment
X12286 N12286 N12287 Segment
X12287 N12287 N12288 Segment
X12288 N12288 N12289 Segment
X12289 N12289 N12290 Segment
X12290 N12290 N12291 Segment
X12291 N12291 N12292 Segment
X12292 N12292 N12293 Segment
X12293 N12293 N12294 Segment
X12294 N12294 N12295 Segment
X12295 N12295 N12296 Segment
X12296 N12296 N12297 Segment
X12297 N12297 N12298 Segment
X12298 N12298 N12299 Segment
X12299 N12299 N12300 Segment
X12300 N12300 N12301 Segment
X12301 N12301 N12302 Segment
X12302 N12302 N12303 Segment
X12303 N12303 N12304 Segment
X12304 N12304 N12305 Segment
X12305 N12305 N12306 Segment
X12306 N12306 N12307 Segment
X12307 N12307 N12308 Segment
X12308 N12308 N12309 Segment
X12309 N12309 N12310 Segment
X12310 N12310 N12311 Segment
X12311 N12311 N12312 Segment
X12312 N12312 N12313 Segment
X12313 N12313 N12314 Segment
X12314 N12314 N12315 Segment
X12315 N12315 N12316 Segment
X12316 N12316 N12317 Segment
X12317 N12317 N12318 Segment
X12318 N12318 N12319 Segment
X12319 N12319 N12320 Segment
X12320 N12320 N12321 Segment
X12321 N12321 N12322 Segment
X12322 N12322 N12323 Segment
X12323 N12323 N12324 Segment
X12324 N12324 N12325 Segment
X12325 N12325 N12326 Segment
X12326 N12326 N12327 Segment
X12327 N12327 N12328 Segment
X12328 N12328 N12329 Segment
X12329 N12329 N12330 Segment
X12330 N12330 N12331 Segment
X12331 N12331 N12332 Segment
X12332 N12332 N12333 Segment
X12333 N12333 N12334 Segment
X12334 N12334 N12335 Segment
X12335 N12335 N12336 Segment
X12336 N12336 N12337 Segment
X12337 N12337 N12338 Segment
X12338 N12338 N12339 Segment
X12339 N12339 N12340 Segment
X12340 N12340 N12341 Segment
X12341 N12341 N12342 Segment
X12342 N12342 N12343 Segment
X12343 N12343 N12344 Segment
X12344 N12344 N12345 Segment
X12345 N12345 N12346 Segment
X12346 N12346 N12347 Segment
X12347 N12347 N12348 Segment
X12348 N12348 N12349 Segment
X12349 N12349 N12350 Segment
X12350 N12350 N12351 Segment
X12351 N12351 N12352 Segment
X12352 N12352 N12353 Segment
X12353 N12353 N12354 Segment
X12354 N12354 N12355 Segment
X12355 N12355 N12356 Segment
X12356 N12356 N12357 Segment
X12357 N12357 N12358 Segment
X12358 N12358 N12359 Segment
X12359 N12359 N12360 Segment
X12360 N12360 N12361 Segment
X12361 N12361 N12362 Segment
X12362 N12362 N12363 Segment
X12363 N12363 N12364 Segment
X12364 N12364 N12365 Segment
X12365 N12365 N12366 Segment
X12366 N12366 N12367 Segment
X12367 N12367 N12368 Segment
X12368 N12368 N12369 Segment
X12369 N12369 N12370 Segment
X12370 N12370 N12371 Segment
X12371 N12371 N12372 Segment
X12372 N12372 N12373 Segment
X12373 N12373 N12374 Segment
X12374 N12374 N12375 Segment
X12375 N12375 N12376 Segment
X12376 N12376 N12377 Segment
X12377 N12377 N12378 Segment
X12378 N12378 N12379 Segment
X12379 N12379 N12380 Segment
X12380 N12380 N12381 Segment
X12381 N12381 N12382 Segment
X12382 N12382 N12383 Segment
X12383 N12383 N12384 Segment
X12384 N12384 N12385 Segment
X12385 N12385 N12386 Segment
X12386 N12386 N12387 Segment
X12387 N12387 N12388 Segment
X12388 N12388 N12389 Segment
X12389 N12389 N12390 Segment
X12390 N12390 N12391 Segment
X12391 N12391 N12392 Segment
X12392 N12392 N12393 Segment
X12393 N12393 N12394 Segment
X12394 N12394 N12395 Segment
X12395 N12395 N12396 Segment
X12396 N12396 N12397 Segment
X12397 N12397 N12398 Segment
X12398 N12398 N12399 Segment
X12399 N12399 N12400 Segment
X12400 N12400 N12401 Segment
X12401 N12401 N12402 Segment
X12402 N12402 N12403 Segment
X12403 N12403 N12404 Segment
X12404 N12404 N12405 Segment
X12405 N12405 N12406 Segment
X12406 N12406 N12407 Segment
X12407 N12407 N12408 Segment
X12408 N12408 N12409 Segment
X12409 N12409 N12410 Segment
X12410 N12410 N12411 Segment
X12411 N12411 N12412 Segment
X12412 N12412 N12413 Segment
X12413 N12413 N12414 Segment
X12414 N12414 N12415 Segment
X12415 N12415 N12416 Segment
X12416 N12416 N12417 Segment
X12417 N12417 N12418 Segment
X12418 N12418 N12419 Segment
X12419 N12419 N12420 Segment
X12420 N12420 N12421 Segment
X12421 N12421 N12422 Segment
X12422 N12422 N12423 Segment
X12423 N12423 N12424 Segment
X12424 N12424 N12425 Segment
X12425 N12425 N12426 Segment
X12426 N12426 N12427 Segment
X12427 N12427 N12428 Segment
X12428 N12428 N12429 Segment
X12429 N12429 N12430 Segment
X12430 N12430 N12431 Segment
X12431 N12431 N12432 Segment
X12432 N12432 N12433 Segment
X12433 N12433 N12434 Segment
X12434 N12434 N12435 Segment
X12435 N12435 N12436 Segment
X12436 N12436 N12437 Segment
X12437 N12437 N12438 Segment
X12438 N12438 N12439 Segment
X12439 N12439 N12440 Segment
X12440 N12440 N12441 Segment
X12441 N12441 N12442 Segment
X12442 N12442 N12443 Segment
X12443 N12443 N12444 Segment
X12444 N12444 N12445 Segment
X12445 N12445 N12446 Segment
X12446 N12446 N12447 Segment
X12447 N12447 N12448 Segment
X12448 N12448 N12449 Segment
X12449 N12449 N12450 Segment
X12450 N12450 N12451 Segment
X12451 N12451 N12452 Segment
X12452 N12452 N12453 Segment
X12453 N12453 N12454 Segment
X12454 N12454 N12455 Segment
X12455 N12455 N12456 Segment
X12456 N12456 N12457 Segment
X12457 N12457 N12458 Segment
X12458 N12458 N12459 Segment
X12459 N12459 N12460 Segment
X12460 N12460 N12461 Segment
X12461 N12461 N12462 Segment
X12462 N12462 N12463 Segment
X12463 N12463 N12464 Segment
X12464 N12464 N12465 Segment
X12465 N12465 N12466 Segment
X12466 N12466 N12467 Segment
X12467 N12467 N12468 Segment
X12468 N12468 N12469 Segment
X12469 N12469 N12470 Segment
X12470 N12470 N12471 Segment
X12471 N12471 N12472 Segment
X12472 N12472 N12473 Segment
X12473 N12473 N12474 Segment
X12474 N12474 N12475 Segment
X12475 N12475 N12476 Segment
X12476 N12476 N12477 Segment
X12477 N12477 N12478 Segment
X12478 N12478 N12479 Segment
X12479 N12479 N12480 Segment
X12480 N12480 N12481 Segment
X12481 N12481 N12482 Segment
X12482 N12482 N12483 Segment
X12483 N12483 N12484 Segment
X12484 N12484 N12485 Segment
X12485 N12485 N12486 Segment
X12486 N12486 N12487 Segment
X12487 N12487 N12488 Segment
X12488 N12488 N12489 Segment
X12489 N12489 N12490 Segment
X12490 N12490 N12491 Segment
X12491 N12491 N12492 Segment
X12492 N12492 N12493 Segment
X12493 N12493 N12494 Segment
X12494 N12494 N12495 Segment
X12495 N12495 N12496 Segment
X12496 N12496 N12497 Segment
X12497 N12497 N12498 Segment
X12498 N12498 N12499 Segment
X12499 N12499 N12500 Segment
X12500 N12500 N12501 Segment
X12501 N12501 N12502 Segment
X12502 N12502 N12503 Segment
X12503 N12503 N12504 Segment
X12504 N12504 N12505 Segment
X12505 N12505 N12506 Segment
X12506 N12506 N12507 Segment
X12507 N12507 N12508 Segment
X12508 N12508 N12509 Segment
X12509 N12509 N12510 Segment
X12510 N12510 N12511 Segment
X12511 N12511 N12512 Segment
X12512 N12512 N12513 Segment
X12513 N12513 N12514 Segment
X12514 N12514 N12515 Segment
X12515 N12515 N12516 Segment
X12516 N12516 N12517 Segment
X12517 N12517 N12518 Segment
X12518 N12518 N12519 Segment
X12519 N12519 N12520 Segment
X12520 N12520 N12521 Segment
X12521 N12521 N12522 Segment
X12522 N12522 N12523 Segment
X12523 N12523 N12524 Segment
X12524 N12524 N12525 Segment
X12525 N12525 N12526 Segment
X12526 N12526 N12527 Segment
X12527 N12527 N12528 Segment
X12528 N12528 N12529 Segment
X12529 N12529 N12530 Segment
X12530 N12530 N12531 Segment
X12531 N12531 N12532 Segment
X12532 N12532 N12533 Segment
X12533 N12533 N12534 Segment
X12534 N12534 N12535 Segment
X12535 N12535 N12536 Segment
X12536 N12536 N12537 Segment
X12537 N12537 N12538 Segment
X12538 N12538 N12539 Segment
X12539 N12539 N12540 Segment
X12540 N12540 N12541 Segment
X12541 N12541 N12542 Segment
X12542 N12542 N12543 Segment
X12543 N12543 N12544 Segment
X12544 N12544 N12545 Segment
X12545 N12545 N12546 Segment
X12546 N12546 N12547 Segment
X12547 N12547 N12548 Segment
X12548 N12548 N12549 Segment
X12549 N12549 N12550 Segment
X12550 N12550 N12551 Segment
X12551 N12551 N12552 Segment
X12552 N12552 N12553 Segment
X12553 N12553 N12554 Segment
X12554 N12554 N12555 Segment
X12555 N12555 N12556 Segment
X12556 N12556 N12557 Segment
X12557 N12557 N12558 Segment
X12558 N12558 N12559 Segment
X12559 N12559 N12560 Segment
X12560 N12560 N12561 Segment
X12561 N12561 N12562 Segment
X12562 N12562 N12563 Segment
X12563 N12563 N12564 Segment
X12564 N12564 N12565 Segment
X12565 N12565 N12566 Segment
X12566 N12566 N12567 Segment
X12567 N12567 N12568 Segment
X12568 N12568 N12569 Segment
X12569 N12569 N12570 Segment
X12570 N12570 N12571 Segment
X12571 N12571 N12572 Segment
X12572 N12572 N12573 Segment
X12573 N12573 N12574 Segment
X12574 N12574 N12575 Segment
X12575 N12575 N12576 Segment
X12576 N12576 N12577 Segment
X12577 N12577 N12578 Segment
X12578 N12578 N12579 Segment
X12579 N12579 N12580 Segment
X12580 N12580 N12581 Segment
X12581 N12581 N12582 Segment
X12582 N12582 N12583 Segment
X12583 N12583 N12584 Segment
X12584 N12584 N12585 Segment
X12585 N12585 N12586 Segment
X12586 N12586 N12587 Segment
X12587 N12587 N12588 Segment
X12588 N12588 N12589 Segment
X12589 N12589 N12590 Segment
X12590 N12590 N12591 Segment
X12591 N12591 N12592 Segment
X12592 N12592 N12593 Segment
X12593 N12593 N12594 Segment
X12594 N12594 N12595 Segment
X12595 N12595 N12596 Segment
X12596 N12596 N12597 Segment
X12597 N12597 N12598 Segment
X12598 N12598 N12599 Segment
X12599 N12599 N12600 Segment
X12600 N12600 N12601 Segment
X12601 N12601 N12602 Segment
X12602 N12602 N12603 Segment
X12603 N12603 N12604 Segment
X12604 N12604 N12605 Segment
X12605 N12605 N12606 Segment
X12606 N12606 N12607 Segment
X12607 N12607 N12608 Segment
X12608 N12608 N12609 Segment
X12609 N12609 N12610 Segment
X12610 N12610 N12611 Segment
X12611 N12611 N12612 Segment
X12612 N12612 N12613 Segment
X12613 N12613 N12614 Segment
X12614 N12614 N12615 Segment
X12615 N12615 N12616 Segment
X12616 N12616 N12617 Segment
X12617 N12617 N12618 Segment
X12618 N12618 N12619 Segment
X12619 N12619 N12620 Segment
X12620 N12620 N12621 Segment
X12621 N12621 N12622 Segment
X12622 N12622 N12623 Segment
X12623 N12623 N12624 Segment
X12624 N12624 N12625 Segment
X12625 N12625 N12626 Segment
X12626 N12626 N12627 Segment
X12627 N12627 N12628 Segment
X12628 N12628 N12629 Segment
X12629 N12629 N12630 Segment
X12630 N12630 N12631 Segment
X12631 N12631 N12632 Segment
X12632 N12632 N12633 Segment
X12633 N12633 N12634 Segment
X12634 N12634 N12635 Segment
X12635 N12635 N12636 Segment
X12636 N12636 N12637 Segment
X12637 N12637 N12638 Segment
X12638 N12638 N12639 Segment
X12639 N12639 N12640 Segment
X12640 N12640 N12641 Segment
X12641 N12641 N12642 Segment
X12642 N12642 N12643 Segment
X12643 N12643 N12644 Segment
X12644 N12644 N12645 Segment
X12645 N12645 N12646 Segment
X12646 N12646 N12647 Segment
X12647 N12647 N12648 Segment
X12648 N12648 N12649 Segment
X12649 N12649 N12650 Segment
X12650 N12650 N12651 Segment
X12651 N12651 N12652 Segment
X12652 N12652 N12653 Segment
X12653 N12653 N12654 Segment
X12654 N12654 N12655 Segment
X12655 N12655 N12656 Segment
X12656 N12656 N12657 Segment
X12657 N12657 N12658 Segment
X12658 N12658 N12659 Segment
X12659 N12659 N12660 Segment
X12660 N12660 N12661 Segment
X12661 N12661 N12662 Segment
X12662 N12662 N12663 Segment
X12663 N12663 N12664 Segment
X12664 N12664 N12665 Segment
X12665 N12665 N12666 Segment
X12666 N12666 N12667 Segment
X12667 N12667 N12668 Segment
X12668 N12668 N12669 Segment
X12669 N12669 N12670 Segment
X12670 N12670 N12671 Segment
X12671 N12671 N12672 Segment
X12672 N12672 N12673 Segment
X12673 N12673 N12674 Segment
X12674 N12674 N12675 Segment
X12675 N12675 N12676 Segment
X12676 N12676 N12677 Segment
X12677 N12677 N12678 Segment
X12678 N12678 N12679 Segment
X12679 N12679 N12680 Segment
X12680 N12680 N12681 Segment
X12681 N12681 N12682 Segment
X12682 N12682 N12683 Segment
X12683 N12683 N12684 Segment
X12684 N12684 N12685 Segment
X12685 N12685 N12686 Segment
X12686 N12686 N12687 Segment
X12687 N12687 N12688 Segment
X12688 N12688 N12689 Segment
X12689 N12689 N12690 Segment
X12690 N12690 N12691 Segment
X12691 N12691 N12692 Segment
X12692 N12692 N12693 Segment
X12693 N12693 N12694 Segment
X12694 N12694 N12695 Segment
X12695 N12695 N12696 Segment
X12696 N12696 N12697 Segment
X12697 N12697 N12698 Segment
X12698 N12698 N12699 Segment
X12699 N12699 N12700 Segment
X12700 N12700 N12701 Segment
X12701 N12701 N12702 Segment
X12702 N12702 N12703 Segment
X12703 N12703 N12704 Segment
X12704 N12704 N12705 Segment
X12705 N12705 N12706 Segment
X12706 N12706 N12707 Segment
X12707 N12707 N12708 Segment
X12708 N12708 N12709 Segment
X12709 N12709 N12710 Segment
X12710 N12710 N12711 Segment
X12711 N12711 N12712 Segment
X12712 N12712 N12713 Segment
X12713 N12713 N12714 Segment
X12714 N12714 N12715 Segment
X12715 N12715 N12716 Segment
X12716 N12716 N12717 Segment
X12717 N12717 N12718 Segment
X12718 N12718 N12719 Segment
X12719 N12719 N12720 Segment
X12720 N12720 N12721 Segment
X12721 N12721 N12722 Segment
X12722 N12722 N12723 Segment
X12723 N12723 N12724 Segment
X12724 N12724 N12725 Segment
X12725 N12725 N12726 Segment
X12726 N12726 N12727 Segment
X12727 N12727 N12728 Segment
X12728 N12728 N12729 Segment
X12729 N12729 N12730 Segment
X12730 N12730 N12731 Segment
X12731 N12731 N12732 Segment
X12732 N12732 N12733 Segment
X12733 N12733 N12734 Segment
X12734 N12734 N12735 Segment
X12735 N12735 N12736 Segment
X12736 N12736 N12737 Segment
X12737 N12737 N12738 Segment
X12738 N12738 N12739 Segment
X12739 N12739 N12740 Segment
X12740 N12740 N12741 Segment
X12741 N12741 N12742 Segment
X12742 N12742 N12743 Segment
X12743 N12743 N12744 Segment
X12744 N12744 N12745 Segment
X12745 N12745 N12746 Segment
X12746 N12746 N12747 Segment
X12747 N12747 N12748 Segment
X12748 N12748 N12749 Segment
X12749 N12749 N12750 Segment
X12750 N12750 N12751 Segment
X12751 N12751 N12752 Segment
X12752 N12752 N12753 Segment
X12753 N12753 N12754 Segment
X12754 N12754 N12755 Segment
X12755 N12755 N12756 Segment
X12756 N12756 N12757 Segment
X12757 N12757 N12758 Segment
X12758 N12758 N12759 Segment
X12759 N12759 N12760 Segment
X12760 N12760 N12761 Segment
X12761 N12761 N12762 Segment
X12762 N12762 N12763 Segment
X12763 N12763 N12764 Segment
X12764 N12764 N12765 Segment
X12765 N12765 N12766 Segment
X12766 N12766 N12767 Segment
X12767 N12767 N12768 Segment
X12768 N12768 N12769 Segment
X12769 N12769 N12770 Segment
X12770 N12770 N12771 Segment
X12771 N12771 N12772 Segment
X12772 N12772 N12773 Segment
X12773 N12773 N12774 Segment
X12774 N12774 N12775 Segment
X12775 N12775 N12776 Segment
X12776 N12776 N12777 Segment
X12777 N12777 N12778 Segment
X12778 N12778 N12779 Segment
X12779 N12779 N12780 Segment
X12780 N12780 N12781 Segment
X12781 N12781 N12782 Segment
X12782 N12782 N12783 Segment
X12783 N12783 N12784 Segment
X12784 N12784 N12785 Segment
X12785 N12785 N12786 Segment
X12786 N12786 N12787 Segment
X12787 N12787 N12788 Segment
X12788 N12788 N12789 Segment
X12789 N12789 N12790 Segment
X12790 N12790 N12791 Segment
X12791 N12791 N12792 Segment
X12792 N12792 N12793 Segment
X12793 N12793 N12794 Segment
X12794 N12794 N12795 Segment
X12795 N12795 N12796 Segment
X12796 N12796 N12797 Segment
X12797 N12797 N12798 Segment
X12798 N12798 N12799 Segment
X12799 N12799 N12800 Segment
X12800 N12800 N12801 Segment
X12801 N12801 N12802 Segment
X12802 N12802 N12803 Segment
X12803 N12803 N12804 Segment
X12804 N12804 N12805 Segment
X12805 N12805 N12806 Segment
X12806 N12806 N12807 Segment
X12807 N12807 N12808 Segment
X12808 N12808 N12809 Segment
X12809 N12809 N12810 Segment
X12810 N12810 N12811 Segment
X12811 N12811 N12812 Segment
X12812 N12812 N12813 Segment
X12813 N12813 N12814 Segment
X12814 N12814 N12815 Segment
X12815 N12815 N12816 Segment
X12816 N12816 N12817 Segment
X12817 N12817 N12818 Segment
X12818 N12818 N12819 Segment
X12819 N12819 N12820 Segment
X12820 N12820 N12821 Segment
X12821 N12821 N12822 Segment
X12822 N12822 N12823 Segment
X12823 N12823 N12824 Segment
X12824 N12824 N12825 Segment
X12825 N12825 N12826 Segment
X12826 N12826 N12827 Segment
X12827 N12827 N12828 Segment
X12828 N12828 N12829 Segment
X12829 N12829 N12830 Segment
X12830 N12830 N12831 Segment
X12831 N12831 N12832 Segment
X12832 N12832 N12833 Segment
X12833 N12833 N12834 Segment
X12834 N12834 N12835 Segment
X12835 N12835 N12836 Segment
X12836 N12836 N12837 Segment
X12837 N12837 N12838 Segment
X12838 N12838 N12839 Segment
X12839 N12839 N12840 Segment
X12840 N12840 N12841 Segment
X12841 N12841 N12842 Segment
X12842 N12842 N12843 Segment
X12843 N12843 N12844 Segment
X12844 N12844 N12845 Segment
X12845 N12845 N12846 Segment
X12846 N12846 N12847 Segment
X12847 N12847 N12848 Segment
X12848 N12848 N12849 Segment
X12849 N12849 N12850 Segment
X12850 N12850 N12851 Segment
X12851 N12851 N12852 Segment
X12852 N12852 N12853 Segment
X12853 N12853 N12854 Segment
X12854 N12854 N12855 Segment
X12855 N12855 N12856 Segment
X12856 N12856 N12857 Segment
X12857 N12857 N12858 Segment
X12858 N12858 N12859 Segment
X12859 N12859 N12860 Segment
X12860 N12860 N12861 Segment
X12861 N12861 N12862 Segment
X12862 N12862 N12863 Segment
X12863 N12863 N12864 Segment
X12864 N12864 N12865 Segment
X12865 N12865 N12866 Segment
X12866 N12866 N12867 Segment
X12867 N12867 N12868 Segment
X12868 N12868 N12869 Segment
X12869 N12869 N12870 Segment
X12870 N12870 N12871 Segment
X12871 N12871 N12872 Segment
X12872 N12872 N12873 Segment
X12873 N12873 N12874 Segment
X12874 N12874 N12875 Segment
X12875 N12875 N12876 Segment
X12876 N12876 N12877 Segment
X12877 N12877 N12878 Segment
X12878 N12878 N12879 Segment
X12879 N12879 N12880 Segment
X12880 N12880 N12881 Segment
X12881 N12881 N12882 Segment
X12882 N12882 N12883 Segment
X12883 N12883 N12884 Segment
X12884 N12884 N12885 Segment
X12885 N12885 N12886 Segment
X12886 N12886 N12887 Segment
X12887 N12887 N12888 Segment
X12888 N12888 N12889 Segment
X12889 N12889 N12890 Segment
X12890 N12890 N12891 Segment
X12891 N12891 N12892 Segment
X12892 N12892 N12893 Segment
X12893 N12893 N12894 Segment
X12894 N12894 N12895 Segment
X12895 N12895 N12896 Segment
X12896 N12896 N12897 Segment
X12897 N12897 N12898 Segment
X12898 N12898 N12899 Segment
X12899 N12899 N12900 Segment
X12900 N12900 N12901 Segment
X12901 N12901 N12902 Segment
X12902 N12902 N12903 Segment
X12903 N12903 N12904 Segment
X12904 N12904 N12905 Segment
X12905 N12905 N12906 Segment
X12906 N12906 N12907 Segment
X12907 N12907 N12908 Segment
X12908 N12908 N12909 Segment
X12909 N12909 N12910 Segment
X12910 N12910 N12911 Segment
X12911 N12911 N12912 Segment
X12912 N12912 N12913 Segment
X12913 N12913 N12914 Segment
X12914 N12914 N12915 Segment
X12915 N12915 N12916 Segment
X12916 N12916 N12917 Segment
X12917 N12917 N12918 Segment
X12918 N12918 N12919 Segment
X12919 N12919 N12920 Segment
X12920 N12920 N12921 Segment
X12921 N12921 N12922 Segment
X12922 N12922 N12923 Segment
X12923 N12923 N12924 Segment
X12924 N12924 N12925 Segment
X12925 N12925 N12926 Segment
X12926 N12926 N12927 Segment
X12927 N12927 N12928 Segment
X12928 N12928 N12929 Segment
X12929 N12929 N12930 Segment
X12930 N12930 N12931 Segment
X12931 N12931 N12932 Segment
X12932 N12932 N12933 Segment
X12933 N12933 N12934 Segment
X12934 N12934 N12935 Segment
X12935 N12935 N12936 Segment
X12936 N12936 N12937 Segment
X12937 N12937 N12938 Segment
X12938 N12938 N12939 Segment
X12939 N12939 N12940 Segment
X12940 N12940 N12941 Segment
X12941 N12941 N12942 Segment
X12942 N12942 N12943 Segment
X12943 N12943 N12944 Segment
X12944 N12944 N12945 Segment
X12945 N12945 N12946 Segment
X12946 N12946 N12947 Segment
X12947 N12947 N12948 Segment
X12948 N12948 N12949 Segment
X12949 N12949 N12950 Segment
X12950 N12950 N12951 Segment
X12951 N12951 N12952 Segment
X12952 N12952 N12953 Segment
X12953 N12953 N12954 Segment
X12954 N12954 N12955 Segment
X12955 N12955 N12956 Segment
X12956 N12956 N12957 Segment
X12957 N12957 N12958 Segment
X12958 N12958 N12959 Segment
X12959 N12959 N12960 Segment
X12960 N12960 N12961 Segment
X12961 N12961 N12962 Segment
X12962 N12962 N12963 Segment
X12963 N12963 N12964 Segment
X12964 N12964 N12965 Segment
X12965 N12965 N12966 Segment
X12966 N12966 N12967 Segment
X12967 N12967 N12968 Segment
X12968 N12968 N12969 Segment
X12969 N12969 N12970 Segment
X12970 N12970 N12971 Segment
X12971 N12971 N12972 Segment
X12972 N12972 N12973 Segment
X12973 N12973 N12974 Segment
X12974 N12974 N12975 Segment
X12975 N12975 N12976 Segment
X12976 N12976 N12977 Segment
X12977 N12977 N12978 Segment
X12978 N12978 N12979 Segment
X12979 N12979 N12980 Segment
X12980 N12980 N12981 Segment
X12981 N12981 N12982 Segment
X12982 N12982 N12983 Segment
X12983 N12983 N12984 Segment
X12984 N12984 N12985 Segment
X12985 N12985 N12986 Segment
X12986 N12986 N12987 Segment
X12987 N12987 N12988 Segment
X12988 N12988 N12989 Segment
X12989 N12989 N12990 Segment
X12990 N12990 N12991 Segment
X12991 N12991 N12992 Segment
X12992 N12992 N12993 Segment
X12993 N12993 N12994 Segment
X12994 N12994 N12995 Segment
X12995 N12995 N12996 Segment
X12996 N12996 N12997 Segment
X12997 N12997 N12998 Segment
X12998 N12998 N12999 Segment
X12999 N12999 N13000 Segment
X13000 N13000 N13001 Segment
X13001 N13001 N13002 Segment
X13002 N13002 N13003 Segment
X13003 N13003 N13004 Segment
X13004 N13004 N13005 Segment
X13005 N13005 N13006 Segment
X13006 N13006 N13007 Segment
X13007 N13007 N13008 Segment
X13008 N13008 N13009 Segment
X13009 N13009 N13010 Segment
X13010 N13010 N13011 Segment
X13011 N13011 N13012 Segment
X13012 N13012 N13013 Segment
X13013 N13013 N13014 Segment
X13014 N13014 N13015 Segment
X13015 N13015 N13016 Segment
X13016 N13016 N13017 Segment
X13017 N13017 N13018 Segment
X13018 N13018 N13019 Segment
X13019 N13019 N13020 Segment
X13020 N13020 N13021 Segment
X13021 N13021 N13022 Segment
X13022 N13022 N13023 Segment
X13023 N13023 N13024 Segment
X13024 N13024 N13025 Segment
X13025 N13025 N13026 Segment
X13026 N13026 N13027 Segment
X13027 N13027 N13028 Segment
X13028 N13028 N13029 Segment
X13029 N13029 N13030 Segment
X13030 N13030 N13031 Segment
X13031 N13031 N13032 Segment
X13032 N13032 N13033 Segment
X13033 N13033 N13034 Segment
X13034 N13034 N13035 Segment
X13035 N13035 N13036 Segment
X13036 N13036 N13037 Segment
X13037 N13037 N13038 Segment
X13038 N13038 N13039 Segment
X13039 N13039 N13040 Segment
X13040 N13040 N13041 Segment
X13041 N13041 N13042 Segment
X13042 N13042 N13043 Segment
X13043 N13043 N13044 Segment
X13044 N13044 N13045 Segment
X13045 N13045 N13046 Segment
X13046 N13046 N13047 Segment
X13047 N13047 N13048 Segment
X13048 N13048 N13049 Segment
X13049 N13049 N13050 Segment
X13050 N13050 N13051 Segment
X13051 N13051 N13052 Segment
X13052 N13052 N13053 Segment
X13053 N13053 N13054 Segment
X13054 N13054 N13055 Segment
X13055 N13055 N13056 Segment
X13056 N13056 N13057 Segment
X13057 N13057 N13058 Segment
X13058 N13058 N13059 Segment
X13059 N13059 N13060 Segment
X13060 N13060 N13061 Segment
X13061 N13061 N13062 Segment
X13062 N13062 N13063 Segment
X13063 N13063 N13064 Segment
X13064 N13064 N13065 Segment
X13065 N13065 N13066 Segment
X13066 N13066 N13067 Segment
X13067 N13067 N13068 Segment
X13068 N13068 N13069 Segment
X13069 N13069 N13070 Segment
X13070 N13070 N13071 Segment
X13071 N13071 N13072 Segment
X13072 N13072 N13073 Segment
X13073 N13073 N13074 Segment
X13074 N13074 N13075 Segment
X13075 N13075 N13076 Segment
X13076 N13076 N13077 Segment
X13077 N13077 N13078 Segment
X13078 N13078 N13079 Segment
X13079 N13079 N13080 Segment
X13080 N13080 N13081 Segment
X13081 N13081 N13082 Segment
X13082 N13082 N13083 Segment
X13083 N13083 N13084 Segment
X13084 N13084 N13085 Segment
X13085 N13085 N13086 Segment
X13086 N13086 N13087 Segment
X13087 N13087 N13088 Segment
X13088 N13088 N13089 Segment
X13089 N13089 N13090 Segment
X13090 N13090 N13091 Segment
X13091 N13091 N13092 Segment
X13092 N13092 N13093 Segment
X13093 N13093 N13094 Segment
X13094 N13094 N13095 Segment
X13095 N13095 N13096 Segment
X13096 N13096 N13097 Segment
X13097 N13097 N13098 Segment
X13098 N13098 N13099 Segment
X13099 N13099 N13100 Segment
X13100 N13100 N13101 Segment
X13101 N13101 N13102 Segment
X13102 N13102 N13103 Segment
X13103 N13103 N13104 Segment
X13104 N13104 N13105 Segment
X13105 N13105 N13106 Segment
X13106 N13106 N13107 Segment
X13107 N13107 N13108 Segment
X13108 N13108 N13109 Segment
X13109 N13109 N13110 Segment
X13110 N13110 N13111 Segment
X13111 N13111 N13112 Segment
X13112 N13112 N13113 Segment
X13113 N13113 N13114 Segment
X13114 N13114 N13115 Segment
X13115 N13115 N13116 Segment
X13116 N13116 N13117 Segment
X13117 N13117 N13118 Segment
X13118 N13118 N13119 Segment
X13119 N13119 N13120 Segment
X13120 N13120 N13121 Segment
X13121 N13121 N13122 Segment
X13122 N13122 N13123 Segment
X13123 N13123 N13124 Segment
X13124 N13124 N13125 Segment
X13125 N13125 N13126 Segment
X13126 N13126 N13127 Segment
X13127 N13127 N13128 Segment
X13128 N13128 N13129 Segment
X13129 N13129 N13130 Segment
X13130 N13130 N13131 Segment
X13131 N13131 N13132 Segment
X13132 N13132 N13133 Segment
X13133 N13133 N13134 Segment
X13134 N13134 N13135 Segment
X13135 N13135 N13136 Segment
X13136 N13136 N13137 Segment
X13137 N13137 N13138 Segment
X13138 N13138 N13139 Segment
X13139 N13139 N13140 Segment
X13140 N13140 N13141 Segment
X13141 N13141 N13142 Segment
X13142 N13142 N13143 Segment
X13143 N13143 N13144 Segment
X13144 N13144 N13145 Segment
X13145 N13145 N13146 Segment
X13146 N13146 N13147 Segment
X13147 N13147 N13148 Segment
X13148 N13148 N13149 Segment
X13149 N13149 N13150 Segment
X13150 N13150 N13151 Segment
X13151 N13151 N13152 Segment
X13152 N13152 N13153 Segment
X13153 N13153 N13154 Segment
X13154 N13154 N13155 Segment
X13155 N13155 N13156 Segment
X13156 N13156 N13157 Segment
X13157 N13157 N13158 Segment
X13158 N13158 N13159 Segment
X13159 N13159 N13160 Segment
X13160 N13160 N13161 Segment
X13161 N13161 N13162 Segment
X13162 N13162 N13163 Segment
X13163 N13163 N13164 Segment
X13164 N13164 N13165 Segment
X13165 N13165 N13166 Segment
X13166 N13166 N13167 Segment
X13167 N13167 N13168 Segment
X13168 N13168 N13169 Segment
X13169 N13169 N13170 Segment
X13170 N13170 N13171 Segment
X13171 N13171 N13172 Segment
X13172 N13172 N13173 Segment
X13173 N13173 N13174 Segment
X13174 N13174 N13175 Segment
X13175 N13175 N13176 Segment
X13176 N13176 N13177 Segment
X13177 N13177 N13178 Segment
X13178 N13178 N13179 Segment
X13179 N13179 N13180 Segment
X13180 N13180 N13181 Segment
X13181 N13181 N13182 Segment
X13182 N13182 N13183 Segment
X13183 N13183 N13184 Segment
X13184 N13184 N13185 Segment
X13185 N13185 N13186 Segment
X13186 N13186 N13187 Segment
X13187 N13187 N13188 Segment
X13188 N13188 N13189 Segment
X13189 N13189 N13190 Segment
X13190 N13190 N13191 Segment
X13191 N13191 N13192 Segment
X13192 N13192 N13193 Segment
X13193 N13193 N13194 Segment
X13194 N13194 N13195 Segment
X13195 N13195 N13196 Segment
X13196 N13196 N13197 Segment
X13197 N13197 N13198 Segment
X13198 N13198 N13199 Segment
X13199 N13199 N13200 Segment
X13200 N13200 N13201 Segment
X13201 N13201 N13202 Segment
X13202 N13202 N13203 Segment
X13203 N13203 N13204 Segment
X13204 N13204 N13205 Segment
X13205 N13205 N13206 Segment
X13206 N13206 N13207 Segment
X13207 N13207 N13208 Segment
X13208 N13208 N13209 Segment
X13209 N13209 N13210 Segment
X13210 N13210 N13211 Segment
X13211 N13211 N13212 Segment
X13212 N13212 N13213 Segment
X13213 N13213 N13214 Segment
X13214 N13214 N13215 Segment
X13215 N13215 N13216 Segment
X13216 N13216 N13217 Segment
X13217 N13217 N13218 Segment
X13218 N13218 N13219 Segment
X13219 N13219 N13220 Segment
X13220 N13220 N13221 Segment
X13221 N13221 N13222 Segment
X13222 N13222 N13223 Segment
X13223 N13223 N13224 Segment
X13224 N13224 N13225 Segment
X13225 N13225 N13226 Segment
X13226 N13226 N13227 Segment
X13227 N13227 N13228 Segment
X13228 N13228 N13229 Segment
X13229 N13229 N13230 Segment
X13230 N13230 N13231 Segment
X13231 N13231 N13232 Segment
X13232 N13232 N13233 Segment
X13233 N13233 N13234 Segment
X13234 N13234 N13235 Segment
X13235 N13235 N13236 Segment
X13236 N13236 N13237 Segment
X13237 N13237 N13238 Segment
X13238 N13238 N13239 Segment
X13239 N13239 N13240 Segment
X13240 N13240 N13241 Segment
X13241 N13241 N13242 Segment
X13242 N13242 N13243 Segment
X13243 N13243 N13244 Segment
X13244 N13244 N13245 Segment
X13245 N13245 N13246 Segment
X13246 N13246 N13247 Segment
X13247 N13247 N13248 Segment
X13248 N13248 N13249 Segment
X13249 N13249 N13250 Segment
X13250 N13250 N13251 Segment
X13251 N13251 N13252 Segment
X13252 N13252 N13253 Segment
X13253 N13253 N13254 Segment
X13254 N13254 N13255 Segment
X13255 N13255 N13256 Segment
X13256 N13256 N13257 Segment
X13257 N13257 N13258 Segment
X13258 N13258 N13259 Segment
X13259 N13259 N13260 Segment
X13260 N13260 N13261 Segment
X13261 N13261 N13262 Segment
X13262 N13262 N13263 Segment
X13263 N13263 N13264 Segment
X13264 N13264 N13265 Segment
X13265 N13265 N13266 Segment
X13266 N13266 N13267 Segment
X13267 N13267 N13268 Segment
X13268 N13268 N13269 Segment
X13269 N13269 N13270 Segment
X13270 N13270 N13271 Segment
X13271 N13271 N13272 Segment
X13272 N13272 N13273 Segment
X13273 N13273 N13274 Segment
X13274 N13274 N13275 Segment
X13275 N13275 N13276 Segment
X13276 N13276 N13277 Segment
X13277 N13277 N13278 Segment
X13278 N13278 N13279 Segment
X13279 N13279 N13280 Segment
X13280 N13280 N13281 Segment
X13281 N13281 N13282 Segment
X13282 N13282 N13283 Segment
X13283 N13283 N13284 Segment
X13284 N13284 N13285 Segment
X13285 N13285 N13286 Segment
X13286 N13286 N13287 Segment
X13287 N13287 N13288 Segment
X13288 N13288 N13289 Segment
X13289 N13289 N13290 Segment
X13290 N13290 N13291 Segment
X13291 N13291 N13292 Segment
X13292 N13292 N13293 Segment
X13293 N13293 N13294 Segment
X13294 N13294 N13295 Segment
X13295 N13295 N13296 Segment
X13296 N13296 N13297 Segment
X13297 N13297 N13298 Segment
X13298 N13298 N13299 Segment
X13299 N13299 N13300 Segment
X13300 N13300 N13301 Segment
X13301 N13301 N13302 Segment
X13302 N13302 N13303 Segment
X13303 N13303 N13304 Segment
X13304 N13304 N13305 Segment
X13305 N13305 N13306 Segment
X13306 N13306 N13307 Segment
X13307 N13307 N13308 Segment
X13308 N13308 N13309 Segment
X13309 N13309 N13310 Segment
X13310 N13310 N13311 Segment
X13311 N13311 N13312 Segment
X13312 N13312 N13313 Segment
X13313 N13313 N13314 Segment
X13314 N13314 N13315 Segment
X13315 N13315 N13316 Segment
X13316 N13316 N13317 Segment
X13317 N13317 N13318 Segment
X13318 N13318 N13319 Segment
X13319 N13319 N13320 Segment
X13320 N13320 N13321 Segment
X13321 N13321 N13322 Segment
X13322 N13322 N13323 Segment
X13323 N13323 N13324 Segment
X13324 N13324 N13325 Segment
X13325 N13325 N13326 Segment
X13326 N13326 N13327 Segment
X13327 N13327 N13328 Segment
X13328 N13328 N13329 Segment
X13329 N13329 N13330 Segment
X13330 N13330 N13331 Segment
X13331 N13331 N13332 Segment
X13332 N13332 N13333 Segment
X13333 N13333 N13334 Segment
X13334 N13334 N13335 Segment
X13335 N13335 N13336 Segment
X13336 N13336 N13337 Segment
X13337 N13337 N13338 Segment
X13338 N13338 N13339 Segment
X13339 N13339 N13340 Segment
X13340 N13340 N13341 Segment
X13341 N13341 N13342 Segment
X13342 N13342 N13343 Segment
X13343 N13343 N13344 Segment
X13344 N13344 N13345 Segment
X13345 N13345 N13346 Segment
X13346 N13346 N13347 Segment
X13347 N13347 N13348 Segment
X13348 N13348 N13349 Segment
X13349 N13349 N13350 Segment
X13350 N13350 N13351 Segment
X13351 N13351 N13352 Segment
X13352 N13352 N13353 Segment
X13353 N13353 N13354 Segment
X13354 N13354 N13355 Segment
X13355 N13355 N13356 Segment
X13356 N13356 N13357 Segment
X13357 N13357 N13358 Segment
X13358 N13358 N13359 Segment
X13359 N13359 N13360 Segment
X13360 N13360 N13361 Segment
X13361 N13361 N13362 Segment
X13362 N13362 N13363 Segment
X13363 N13363 N13364 Segment
X13364 N13364 N13365 Segment
X13365 N13365 N13366 Segment
X13366 N13366 N13367 Segment
X13367 N13367 N13368 Segment
X13368 N13368 N13369 Segment
X13369 N13369 N13370 Segment
X13370 N13370 N13371 Segment
X13371 N13371 N13372 Segment
X13372 N13372 N13373 Segment
X13373 N13373 N13374 Segment
X13374 N13374 N13375 Segment
X13375 N13375 N13376 Segment
X13376 N13376 N13377 Segment
X13377 N13377 N13378 Segment
X13378 N13378 N13379 Segment
X13379 N13379 N13380 Segment
X13380 N13380 N13381 Segment
X13381 N13381 N13382 Segment
X13382 N13382 N13383 Segment
X13383 N13383 N13384 Segment
X13384 N13384 N13385 Segment
X13385 N13385 N13386 Segment
X13386 N13386 N13387 Segment
X13387 N13387 N13388 Segment
X13388 N13388 N13389 Segment
X13389 N13389 N13390 Segment
X13390 N13390 N13391 Segment
X13391 N13391 N13392 Segment
X13392 N13392 N13393 Segment
X13393 N13393 N13394 Segment
X13394 N13394 N13395 Segment
X13395 N13395 N13396 Segment
X13396 N13396 N13397 Segment
X13397 N13397 N13398 Segment
X13398 N13398 N13399 Segment
X13399 N13399 N13400 Segment
X13400 N13400 N13401 Segment
X13401 N13401 N13402 Segment
X13402 N13402 N13403 Segment
X13403 N13403 N13404 Segment
X13404 N13404 N13405 Segment
X13405 N13405 N13406 Segment
X13406 N13406 N13407 Segment
X13407 N13407 N13408 Segment
X13408 N13408 N13409 Segment
X13409 N13409 N13410 Segment
X13410 N13410 N13411 Segment
X13411 N13411 N13412 Segment
X13412 N13412 N13413 Segment
X13413 N13413 N13414 Segment
X13414 N13414 N13415 Segment
X13415 N13415 N13416 Segment
X13416 N13416 N13417 Segment
X13417 N13417 N13418 Segment
X13418 N13418 N13419 Segment
X13419 N13419 N13420 Segment
X13420 N13420 N13421 Segment
X13421 N13421 N13422 Segment
X13422 N13422 N13423 Segment
X13423 N13423 N13424 Segment
X13424 N13424 N13425 Segment
X13425 N13425 N13426 Segment
X13426 N13426 N13427 Segment
X13427 N13427 N13428 Segment
X13428 N13428 N13429 Segment
X13429 N13429 N13430 Segment
X13430 N13430 N13431 Segment
X13431 N13431 N13432 Segment
X13432 N13432 N13433 Segment
X13433 N13433 N13434 Segment
X13434 N13434 N13435 Segment
X13435 N13435 N13436 Segment
X13436 N13436 N13437 Segment
X13437 N13437 N13438 Segment
X13438 N13438 N13439 Segment
X13439 N13439 N13440 Segment
X13440 N13440 N13441 Segment
X13441 N13441 N13442 Segment
X13442 N13442 N13443 Segment
X13443 N13443 N13444 Segment
X13444 N13444 N13445 Segment
X13445 N13445 N13446 Segment
X13446 N13446 N13447 Segment
X13447 N13447 N13448 Segment
X13448 N13448 N13449 Segment
X13449 N13449 N13450 Segment
X13450 N13450 N13451 Segment
X13451 N13451 N13452 Segment
X13452 N13452 N13453 Segment
X13453 N13453 N13454 Segment
X13454 N13454 N13455 Segment
X13455 N13455 N13456 Segment
X13456 N13456 N13457 Segment
X13457 N13457 N13458 Segment
X13458 N13458 N13459 Segment
X13459 N13459 N13460 Segment
X13460 N13460 N13461 Segment
X13461 N13461 N13462 Segment
X13462 N13462 N13463 Segment
X13463 N13463 N13464 Segment
X13464 N13464 N13465 Segment
X13465 N13465 N13466 Segment
X13466 N13466 N13467 Segment
X13467 N13467 N13468 Segment
X13468 N13468 N13469 Segment
X13469 N13469 N13470 Segment
X13470 N13470 N13471 Segment
X13471 N13471 N13472 Segment
X13472 N13472 N13473 Segment
X13473 N13473 N13474 Segment
X13474 N13474 N13475 Segment
X13475 N13475 N13476 Segment
X13476 N13476 N13477 Segment
X13477 N13477 N13478 Segment
X13478 N13478 N13479 Segment
X13479 N13479 N13480 Segment
X13480 N13480 N13481 Segment
X13481 N13481 N13482 Segment
X13482 N13482 N13483 Segment
X13483 N13483 N13484 Segment
X13484 N13484 N13485 Segment
X13485 N13485 N13486 Segment
X13486 N13486 N13487 Segment
X13487 N13487 N13488 Segment
X13488 N13488 N13489 Segment
X13489 N13489 N13490 Segment
X13490 N13490 N13491 Segment
X13491 N13491 N13492 Segment
X13492 N13492 N13493 Segment
X13493 N13493 N13494 Segment
X13494 N13494 N13495 Segment
X13495 N13495 N13496 Segment
X13496 N13496 N13497 Segment
X13497 N13497 N13498 Segment
X13498 N13498 N13499 Segment
X13499 N13499 N13500 Segment
X13500 N13500 N13501 Segment
X13501 N13501 N13502 Segment
X13502 N13502 N13503 Segment
X13503 N13503 N13504 Segment
X13504 N13504 N13505 Segment
X13505 N13505 N13506 Segment
X13506 N13506 N13507 Segment
X13507 N13507 N13508 Segment
X13508 N13508 N13509 Segment
X13509 N13509 N13510 Segment
X13510 N13510 N13511 Segment
X13511 N13511 N13512 Segment
X13512 N13512 N13513 Segment
X13513 N13513 N13514 Segment
X13514 N13514 N13515 Segment
X13515 N13515 N13516 Segment
X13516 N13516 N13517 Segment
X13517 N13517 N13518 Segment
X13518 N13518 N13519 Segment
X13519 N13519 N13520 Segment
X13520 N13520 N13521 Segment
X13521 N13521 N13522 Segment
X13522 N13522 N13523 Segment
X13523 N13523 N13524 Segment
X13524 N13524 N13525 Segment
X13525 N13525 N13526 Segment
X13526 N13526 N13527 Segment
X13527 N13527 N13528 Segment
X13528 N13528 N13529 Segment
X13529 N13529 N13530 Segment
X13530 N13530 N13531 Segment
X13531 N13531 N13532 Segment
X13532 N13532 N13533 Segment
X13533 N13533 N13534 Segment
X13534 N13534 N13535 Segment
X13535 N13535 N13536 Segment
X13536 N13536 N13537 Segment
X13537 N13537 N13538 Segment
X13538 N13538 N13539 Segment
X13539 N13539 N13540 Segment
X13540 N13540 N13541 Segment
X13541 N13541 N13542 Segment
X13542 N13542 N13543 Segment
X13543 N13543 N13544 Segment
X13544 N13544 N13545 Segment
X13545 N13545 N13546 Segment
X13546 N13546 N13547 Segment
X13547 N13547 N13548 Segment
X13548 N13548 N13549 Segment
X13549 N13549 N13550 Segment
X13550 N13550 N13551 Segment
X13551 N13551 N13552 Segment
X13552 N13552 N13553 Segment
X13553 N13553 N13554 Segment
X13554 N13554 N13555 Segment
X13555 N13555 N13556 Segment
X13556 N13556 N13557 Segment
X13557 N13557 N13558 Segment
X13558 N13558 N13559 Segment
X13559 N13559 N13560 Segment
X13560 N13560 N13561 Segment
X13561 N13561 N13562 Segment
X13562 N13562 N13563 Segment
X13563 N13563 N13564 Segment
X13564 N13564 N13565 Segment
X13565 N13565 N13566 Segment
X13566 N13566 N13567 Segment
X13567 N13567 N13568 Segment
X13568 N13568 N13569 Segment
X13569 N13569 N13570 Segment
X13570 N13570 N13571 Segment
X13571 N13571 N13572 Segment
X13572 N13572 N13573 Segment
X13573 N13573 N13574 Segment
X13574 N13574 N13575 Segment
X13575 N13575 N13576 Segment
X13576 N13576 N13577 Segment
X13577 N13577 N13578 Segment
X13578 N13578 N13579 Segment
X13579 N13579 N13580 Segment
X13580 N13580 N13581 Segment
X13581 N13581 N13582 Segment
X13582 N13582 N13583 Segment
X13583 N13583 N13584 Segment
X13584 N13584 N13585 Segment
X13585 N13585 N13586 Segment
X13586 N13586 N13587 Segment
X13587 N13587 N13588 Segment
X13588 N13588 N13589 Segment
X13589 N13589 N13590 Segment
X13590 N13590 N13591 Segment
X13591 N13591 N13592 Segment
X13592 N13592 N13593 Segment
X13593 N13593 N13594 Segment
X13594 N13594 N13595 Segment
X13595 N13595 N13596 Segment
X13596 N13596 N13597 Segment
X13597 N13597 N13598 Segment
X13598 N13598 N13599 Segment
X13599 N13599 N13600 Segment
X13600 N13600 N13601 Segment
X13601 N13601 N13602 Segment
X13602 N13602 N13603 Segment
X13603 N13603 N13604 Segment
X13604 N13604 N13605 Segment
X13605 N13605 N13606 Segment
X13606 N13606 N13607 Segment
X13607 N13607 N13608 Segment
X13608 N13608 N13609 Segment
X13609 N13609 N13610 Segment
X13610 N13610 N13611 Segment
X13611 N13611 N13612 Segment
X13612 N13612 N13613 Segment
X13613 N13613 N13614 Segment
X13614 N13614 N13615 Segment
X13615 N13615 N13616 Segment
X13616 N13616 N13617 Segment
X13617 N13617 N13618 Segment
X13618 N13618 N13619 Segment
X13619 N13619 N13620 Segment
X13620 N13620 N13621 Segment
X13621 N13621 N13622 Segment
X13622 N13622 N13623 Segment
X13623 N13623 N13624 Segment
X13624 N13624 N13625 Segment
X13625 N13625 N13626 Segment
X13626 N13626 N13627 Segment
X13627 N13627 N13628 Segment
X13628 N13628 N13629 Segment
X13629 N13629 N13630 Segment
X13630 N13630 N13631 Segment
X13631 N13631 N13632 Segment
X13632 N13632 N13633 Segment
X13633 N13633 N13634 Segment
X13634 N13634 N13635 Segment
X13635 N13635 N13636 Segment
X13636 N13636 N13637 Segment
X13637 N13637 N13638 Segment
X13638 N13638 N13639 Segment
X13639 N13639 N13640 Segment
X13640 N13640 N13641 Segment
X13641 N13641 N13642 Segment
X13642 N13642 N13643 Segment
X13643 N13643 N13644 Segment
X13644 N13644 N13645 Segment
X13645 N13645 N13646 Segment
X13646 N13646 N13647 Segment
X13647 N13647 N13648 Segment
X13648 N13648 N13649 Segment
X13649 N13649 N13650 Segment
X13650 N13650 N13651 Segment
X13651 N13651 N13652 Segment
X13652 N13652 N13653 Segment
X13653 N13653 N13654 Segment
X13654 N13654 N13655 Segment
X13655 N13655 N13656 Segment
X13656 N13656 N13657 Segment
X13657 N13657 N13658 Segment
X13658 N13658 N13659 Segment
X13659 N13659 N13660 Segment
X13660 N13660 N13661 Segment
X13661 N13661 N13662 Segment
X13662 N13662 N13663 Segment
X13663 N13663 N13664 Segment
X13664 N13664 N13665 Segment
X13665 N13665 N13666 Segment
X13666 N13666 N13667 Segment
X13667 N13667 N13668 Segment
X13668 N13668 N13669 Segment
X13669 N13669 N13670 Segment
X13670 N13670 N13671 Segment
X13671 N13671 N13672 Segment
X13672 N13672 N13673 Segment
X13673 N13673 N13674 Segment
X13674 N13674 N13675 Segment
X13675 N13675 N13676 Segment
X13676 N13676 N13677 Segment
X13677 N13677 N13678 Segment
X13678 N13678 N13679 Segment
X13679 N13679 N13680 Segment
X13680 N13680 N13681 Segment
X13681 N13681 N13682 Segment
X13682 N13682 N13683 Segment
X13683 N13683 N13684 Segment
X13684 N13684 N13685 Segment
X13685 N13685 N13686 Segment
X13686 N13686 N13687 Segment
X13687 N13687 N13688 Segment
X13688 N13688 N13689 Segment
X13689 N13689 N13690 Segment
X13690 N13690 N13691 Segment
X13691 N13691 N13692 Segment
X13692 N13692 N13693 Segment
X13693 N13693 N13694 Segment
X13694 N13694 N13695 Segment
X13695 N13695 N13696 Segment
X13696 N13696 N13697 Segment
X13697 N13697 N13698 Segment
X13698 N13698 N13699 Segment
X13699 N13699 N13700 Segment
X13700 N13700 N13701 Segment
X13701 N13701 N13702 Segment
X13702 N13702 N13703 Segment
X13703 N13703 N13704 Segment
X13704 N13704 N13705 Segment
X13705 N13705 N13706 Segment
X13706 N13706 N13707 Segment
X13707 N13707 N13708 Segment
X13708 N13708 N13709 Segment
X13709 N13709 N13710 Segment
X13710 N13710 N13711 Segment
X13711 N13711 N13712 Segment
X13712 N13712 N13713 Segment
X13713 N13713 N13714 Segment
X13714 N13714 N13715 Segment
X13715 N13715 N13716 Segment
X13716 N13716 N13717 Segment
X13717 N13717 N13718 Segment
X13718 N13718 N13719 Segment
X13719 N13719 N13720 Segment
X13720 N13720 N13721 Segment
X13721 N13721 N13722 Segment
X13722 N13722 N13723 Segment
X13723 N13723 N13724 Segment
X13724 N13724 N13725 Segment
X13725 N13725 N13726 Segment
X13726 N13726 N13727 Segment
X13727 N13727 N13728 Segment
X13728 N13728 N13729 Segment
X13729 N13729 N13730 Segment
X13730 N13730 N13731 Segment
X13731 N13731 N13732 Segment
X13732 N13732 N13733 Segment
X13733 N13733 N13734 Segment
X13734 N13734 N13735 Segment
X13735 N13735 N13736 Segment
X13736 N13736 N13737 Segment
X13737 N13737 N13738 Segment
X13738 N13738 N13739 Segment
X13739 N13739 N13740 Segment
X13740 N13740 N13741 Segment
X13741 N13741 N13742 Segment
X13742 N13742 N13743 Segment
X13743 N13743 N13744 Segment
X13744 N13744 N13745 Segment
X13745 N13745 N13746 Segment
X13746 N13746 N13747 Segment
X13747 N13747 N13748 Segment
X13748 N13748 N13749 Segment
X13749 N13749 N13750 Segment
X13750 N13750 N13751 Segment
X13751 N13751 N13752 Segment
X13752 N13752 N13753 Segment
X13753 N13753 N13754 Segment
X13754 N13754 N13755 Segment
X13755 N13755 N13756 Segment
X13756 N13756 N13757 Segment
X13757 N13757 N13758 Segment
X13758 N13758 N13759 Segment
X13759 N13759 N13760 Segment
X13760 N13760 N13761 Segment
X13761 N13761 N13762 Segment
X13762 N13762 N13763 Segment
X13763 N13763 N13764 Segment
X13764 N13764 N13765 Segment
X13765 N13765 N13766 Segment
X13766 N13766 N13767 Segment
X13767 N13767 N13768 Segment
X13768 N13768 N13769 Segment
X13769 N13769 N13770 Segment
X13770 N13770 N13771 Segment
X13771 N13771 N13772 Segment
X13772 N13772 N13773 Segment
X13773 N13773 N13774 Segment
X13774 N13774 N13775 Segment
X13775 N13775 N13776 Segment
X13776 N13776 N13777 Segment
X13777 N13777 N13778 Segment
X13778 N13778 N13779 Segment
X13779 N13779 N13780 Segment
X13780 N13780 N13781 Segment
X13781 N13781 N13782 Segment
X13782 N13782 N13783 Segment
X13783 N13783 N13784 Segment
X13784 N13784 N13785 Segment
X13785 N13785 N13786 Segment
X13786 N13786 N13787 Segment
X13787 N13787 N13788 Segment
X13788 N13788 N13789 Segment
X13789 N13789 N13790 Segment
X13790 N13790 N13791 Segment
X13791 N13791 N13792 Segment
X13792 N13792 N13793 Segment
X13793 N13793 N13794 Segment
X13794 N13794 N13795 Segment
X13795 N13795 N13796 Segment
X13796 N13796 N13797 Segment
X13797 N13797 N13798 Segment
X13798 N13798 N13799 Segment
X13799 N13799 N13800 Segment
X13800 N13800 N13801 Segment
X13801 N13801 N13802 Segment
X13802 N13802 N13803 Segment
X13803 N13803 N13804 Segment
X13804 N13804 N13805 Segment
X13805 N13805 N13806 Segment
X13806 N13806 N13807 Segment
X13807 N13807 N13808 Segment
X13808 N13808 N13809 Segment
X13809 N13809 N13810 Segment
X13810 N13810 N13811 Segment
X13811 N13811 N13812 Segment
X13812 N13812 N13813 Segment
X13813 N13813 N13814 Segment
X13814 N13814 N13815 Segment
X13815 N13815 N13816 Segment
X13816 N13816 N13817 Segment
X13817 N13817 N13818 Segment
X13818 N13818 N13819 Segment
X13819 N13819 N13820 Segment
X13820 N13820 N13821 Segment
X13821 N13821 N13822 Segment
X13822 N13822 N13823 Segment
X13823 N13823 N13824 Segment
X13824 N13824 N13825 Segment
X13825 N13825 N13826 Segment
X13826 N13826 N13827 Segment
X13827 N13827 N13828 Segment
X13828 N13828 N13829 Segment
X13829 N13829 N13830 Segment
X13830 N13830 N13831 Segment
X13831 N13831 N13832 Segment
X13832 N13832 N13833 Segment
X13833 N13833 N13834 Segment
X13834 N13834 N13835 Segment
X13835 N13835 N13836 Segment
X13836 N13836 N13837 Segment
X13837 N13837 N13838 Segment
X13838 N13838 N13839 Segment
X13839 N13839 N13840 Segment
X13840 N13840 N13841 Segment
X13841 N13841 N13842 Segment
X13842 N13842 N13843 Segment
X13843 N13843 N13844 Segment
X13844 N13844 N13845 Segment
X13845 N13845 N13846 Segment
X13846 N13846 N13847 Segment
X13847 N13847 N13848 Segment
X13848 N13848 N13849 Segment
X13849 N13849 N13850 Segment
X13850 N13850 N13851 Segment
X13851 N13851 N13852 Segment
X13852 N13852 N13853 Segment
X13853 N13853 N13854 Segment
X13854 N13854 N13855 Segment
X13855 N13855 N13856 Segment
X13856 N13856 N13857 Segment
X13857 N13857 N13858 Segment
X13858 N13858 N13859 Segment
X13859 N13859 N13860 Segment
X13860 N13860 N13861 Segment
X13861 N13861 N13862 Segment
X13862 N13862 N13863 Segment
X13863 N13863 N13864 Segment
X13864 N13864 N13865 Segment
X13865 N13865 N13866 Segment
X13866 N13866 N13867 Segment
X13867 N13867 N13868 Segment
X13868 N13868 N13869 Segment
X13869 N13869 N13870 Segment
X13870 N13870 N13871 Segment
X13871 N13871 N13872 Segment
X13872 N13872 N13873 Segment
X13873 N13873 N13874 Segment
X13874 N13874 N13875 Segment
X13875 N13875 N13876 Segment
X13876 N13876 N13877 Segment
X13877 N13877 N13878 Segment
X13878 N13878 N13879 Segment
X13879 N13879 N13880 Segment
X13880 N13880 N13881 Segment
X13881 N13881 N13882 Segment
X13882 N13882 N13883 Segment
X13883 N13883 N13884 Segment
X13884 N13884 N13885 Segment
X13885 N13885 N13886 Segment
X13886 N13886 N13887 Segment
X13887 N13887 N13888 Segment
X13888 N13888 N13889 Segment
X13889 N13889 N13890 Segment
X13890 N13890 N13891 Segment
X13891 N13891 N13892 Segment
X13892 N13892 N13893 Segment
X13893 N13893 N13894 Segment
X13894 N13894 N13895 Segment
X13895 N13895 N13896 Segment
X13896 N13896 N13897 Segment
X13897 N13897 N13898 Segment
X13898 N13898 N13899 Segment
X13899 N13899 N13900 Segment
X13900 N13900 N13901 Segment
X13901 N13901 N13902 Segment
X13902 N13902 N13903 Segment
X13903 N13903 N13904 Segment
X13904 N13904 N13905 Segment
X13905 N13905 N13906 Segment
X13906 N13906 N13907 Segment
X13907 N13907 N13908 Segment
X13908 N13908 N13909 Segment
X13909 N13909 N13910 Segment
X13910 N13910 N13911 Segment
X13911 N13911 N13912 Segment
X13912 N13912 N13913 Segment
X13913 N13913 N13914 Segment
X13914 N13914 N13915 Segment
X13915 N13915 N13916 Segment
X13916 N13916 N13917 Segment
X13917 N13917 N13918 Segment
X13918 N13918 N13919 Segment
X13919 N13919 N13920 Segment
X13920 N13920 N13921 Segment
X13921 N13921 N13922 Segment
X13922 N13922 N13923 Segment
X13923 N13923 N13924 Segment
X13924 N13924 N13925 Segment
X13925 N13925 N13926 Segment
X13926 N13926 N13927 Segment
X13927 N13927 N13928 Segment
X13928 N13928 N13929 Segment
X13929 N13929 N13930 Segment
X13930 N13930 N13931 Segment
X13931 N13931 N13932 Segment
X13932 N13932 N13933 Segment
X13933 N13933 N13934 Segment
X13934 N13934 N13935 Segment
X13935 N13935 N13936 Segment
X13936 N13936 N13937 Segment
X13937 N13937 N13938 Segment
X13938 N13938 N13939 Segment
X13939 N13939 N13940 Segment
X13940 N13940 N13941 Segment
X13941 N13941 N13942 Segment
X13942 N13942 N13943 Segment
X13943 N13943 N13944 Segment
X13944 N13944 N13945 Segment
X13945 N13945 N13946 Segment
X13946 N13946 N13947 Segment
X13947 N13947 N13948 Segment
X13948 N13948 N13949 Segment
X13949 N13949 N13950 Segment
X13950 N13950 N13951 Segment
X13951 N13951 N13952 Segment
X13952 N13952 N13953 Segment
X13953 N13953 N13954 Segment
X13954 N13954 N13955 Segment
X13955 N13955 N13956 Segment
X13956 N13956 N13957 Segment
X13957 N13957 N13958 Segment
X13958 N13958 N13959 Segment
X13959 N13959 N13960 Segment
X13960 N13960 N13961 Segment
X13961 N13961 N13962 Segment
X13962 N13962 N13963 Segment
X13963 N13963 N13964 Segment
X13964 N13964 N13965 Segment
X13965 N13965 N13966 Segment
X13966 N13966 N13967 Segment
X13967 N13967 N13968 Segment
X13968 N13968 N13969 Segment
X13969 N13969 N13970 Segment
X13970 N13970 N13971 Segment
X13971 N13971 N13972 Segment
X13972 N13972 N13973 Segment
X13973 N13973 N13974 Segment
X13974 N13974 N13975 Segment
X13975 N13975 N13976 Segment
X13976 N13976 N13977 Segment
X13977 N13977 N13978 Segment
X13978 N13978 N13979 Segment
X13979 N13979 N13980 Segment
X13980 N13980 N13981 Segment
X13981 N13981 N13982 Segment
X13982 N13982 N13983 Segment
X13983 N13983 N13984 Segment
X13984 N13984 N13985 Segment
X13985 N13985 N13986 Segment
X13986 N13986 N13987 Segment
X13987 N13987 N13988 Segment
X13988 N13988 N13989 Segment
X13989 N13989 N13990 Segment
X13990 N13990 N13991 Segment
X13991 N13991 N13992 Segment
X13992 N13992 N13993 Segment
X13993 N13993 N13994 Segment
X13994 N13994 N13995 Segment
X13995 N13995 N13996 Segment
X13996 N13996 N13997 Segment
X13997 N13997 N13998 Segment
X13998 N13998 N13999 Segment
X13999 N13999 N14000 Segment
X14000 N14000 N14001 Segment
X14001 N14001 N14002 Segment
X14002 N14002 N14003 Segment
X14003 N14003 N14004 Segment
X14004 N14004 N14005 Segment
X14005 N14005 N14006 Segment
X14006 N14006 N14007 Segment
X14007 N14007 N14008 Segment
X14008 N14008 N14009 Segment
X14009 N14009 N14010 Segment
X14010 N14010 N14011 Segment
X14011 N14011 N14012 Segment
X14012 N14012 N14013 Segment
X14013 N14013 N14014 Segment
X14014 N14014 N14015 Segment
X14015 N14015 N14016 Segment
X14016 N14016 N14017 Segment
X14017 N14017 N14018 Segment
X14018 N14018 N14019 Segment
X14019 N14019 N14020 Segment
X14020 N14020 N14021 Segment
X14021 N14021 N14022 Segment
X14022 N14022 N14023 Segment
X14023 N14023 N14024 Segment
X14024 N14024 N14025 Segment
X14025 N14025 N14026 Segment
X14026 N14026 N14027 Segment
X14027 N14027 N14028 Segment
X14028 N14028 N14029 Segment
X14029 N14029 N14030 Segment
X14030 N14030 N14031 Segment
X14031 N14031 N14032 Segment
X14032 N14032 N14033 Segment
X14033 N14033 N14034 Segment
X14034 N14034 N14035 Segment
X14035 N14035 N14036 Segment
X14036 N14036 N14037 Segment
X14037 N14037 N14038 Segment
X14038 N14038 N14039 Segment
X14039 N14039 N14040 Segment
X14040 N14040 N14041 Segment
X14041 N14041 N14042 Segment
X14042 N14042 N14043 Segment
X14043 N14043 N14044 Segment
X14044 N14044 N14045 Segment
X14045 N14045 N14046 Segment
X14046 N14046 N14047 Segment
X14047 N14047 N14048 Segment
X14048 N14048 N14049 Segment
X14049 N14049 N14050 Segment
X14050 N14050 N14051 Segment
X14051 N14051 N14052 Segment
X14052 N14052 N14053 Segment
X14053 N14053 N14054 Segment
X14054 N14054 N14055 Segment
X14055 N14055 N14056 Segment
X14056 N14056 N14057 Segment
X14057 N14057 N14058 Segment
X14058 N14058 N14059 Segment
X14059 N14059 N14060 Segment
X14060 N14060 N14061 Segment
X14061 N14061 N14062 Segment
X14062 N14062 N14063 Segment
X14063 N14063 N14064 Segment
X14064 N14064 N14065 Segment
X14065 N14065 N14066 Segment
X14066 N14066 N14067 Segment
X14067 N14067 N14068 Segment
X14068 N14068 N14069 Segment
X14069 N14069 N14070 Segment
X14070 N14070 N14071 Segment
X14071 N14071 N14072 Segment
X14072 N14072 N14073 Segment
X14073 N14073 N14074 Segment
X14074 N14074 N14075 Segment
X14075 N14075 N14076 Segment
X14076 N14076 N14077 Segment
X14077 N14077 N14078 Segment
X14078 N14078 N14079 Segment
X14079 N14079 N14080 Segment
X14080 N14080 N14081 Segment
X14081 N14081 N14082 Segment
X14082 N14082 N14083 Segment
X14083 N14083 N14084 Segment
X14084 N14084 N14085 Segment
X14085 N14085 N14086 Segment
X14086 N14086 N14087 Segment
X14087 N14087 N14088 Segment
X14088 N14088 N14089 Segment
X14089 N14089 N14090 Segment
X14090 N14090 N14091 Segment
X14091 N14091 N14092 Segment
X14092 N14092 N14093 Segment
X14093 N14093 N14094 Segment
X14094 N14094 N14095 Segment
X14095 N14095 N14096 Segment
X14096 N14096 N14097 Segment
X14097 N14097 N14098 Segment
X14098 N14098 N14099 Segment
X14099 N14099 N14100 Segment
X14100 N14100 N14101 Segment
X14101 N14101 N14102 Segment
X14102 N14102 N14103 Segment
X14103 N14103 N14104 Segment
X14104 N14104 N14105 Segment
X14105 N14105 N14106 Segment
X14106 N14106 N14107 Segment
X14107 N14107 N14108 Segment
X14108 N14108 N14109 Segment
X14109 N14109 N14110 Segment
X14110 N14110 N14111 Segment
X14111 N14111 N14112 Segment
X14112 N14112 N14113 Segment
X14113 N14113 N14114 Segment
X14114 N14114 N14115 Segment
X14115 N14115 N14116 Segment
X14116 N14116 N14117 Segment
X14117 N14117 N14118 Segment
X14118 N14118 N14119 Segment
X14119 N14119 N14120 Segment
X14120 N14120 N14121 Segment
X14121 N14121 N14122 Segment
X14122 N14122 N14123 Segment
X14123 N14123 N14124 Segment
X14124 N14124 N14125 Segment
X14125 N14125 N14126 Segment
X14126 N14126 N14127 Segment
X14127 N14127 N14128 Segment
X14128 N14128 N14129 Segment
X14129 N14129 N14130 Segment
X14130 N14130 N14131 Segment
X14131 N14131 N14132 Segment
X14132 N14132 N14133 Segment
X14133 N14133 N14134 Segment
X14134 N14134 N14135 Segment
X14135 N14135 N14136 Segment
X14136 N14136 N14137 Segment
X14137 N14137 N14138 Segment
X14138 N14138 N14139 Segment
X14139 N14139 N14140 Segment
X14140 N14140 N14141 Segment
X14141 N14141 N14142 Segment
X14142 N14142 N14143 Segment
X14143 N14143 N14144 Segment
X14144 N14144 N14145 Segment
X14145 N14145 N14146 Segment
X14146 N14146 N14147 Segment
X14147 N14147 N14148 Segment
X14148 N14148 N14149 Segment
X14149 N14149 N14150 Segment
X14150 N14150 N14151 Segment
X14151 N14151 N14152 Segment
X14152 N14152 N14153 Segment
X14153 N14153 N14154 Segment
X14154 N14154 N14155 Segment
X14155 N14155 N14156 Segment
X14156 N14156 N14157 Segment
X14157 N14157 N14158 Segment
X14158 N14158 N14159 Segment
X14159 N14159 N14160 Segment
X14160 N14160 N14161 Segment
X14161 N14161 N14162 Segment
X14162 N14162 N14163 Segment
X14163 N14163 N14164 Segment
X14164 N14164 N14165 Segment
X14165 N14165 N14166 Segment
X14166 N14166 N14167 Segment
X14167 N14167 N14168 Segment
X14168 N14168 N14169 Segment
X14169 N14169 N14170 Segment
X14170 N14170 N14171 Segment
X14171 N14171 N14172 Segment
X14172 N14172 N14173 Segment
X14173 N14173 N14174 Segment
X14174 N14174 N14175 Segment
X14175 N14175 N14176 Segment
X14176 N14176 N14177 Segment
X14177 N14177 N14178 Segment
X14178 N14178 N14179 Segment
X14179 N14179 N14180 Segment
X14180 N14180 N14181 Segment
X14181 N14181 N14182 Segment
X14182 N14182 N14183 Segment
X14183 N14183 N14184 Segment
X14184 N14184 N14185 Segment
X14185 N14185 N14186 Segment
X14186 N14186 N14187 Segment
X14187 N14187 N14188 Segment
X14188 N14188 N14189 Segment
X14189 N14189 N14190 Segment
X14190 N14190 N14191 Segment
X14191 N14191 N14192 Segment
X14192 N14192 N14193 Segment
X14193 N14193 N14194 Segment
X14194 N14194 N14195 Segment
X14195 N14195 N14196 Segment
X14196 N14196 N14197 Segment
X14197 N14197 N14198 Segment
X14198 N14198 N14199 Segment
X14199 N14199 N14200 Segment
X14200 N14200 N14201 Segment
X14201 N14201 N14202 Segment
X14202 N14202 N14203 Segment
X14203 N14203 N14204 Segment
X14204 N14204 N14205 Segment
X14205 N14205 N14206 Segment
X14206 N14206 N14207 Segment
X14207 N14207 N14208 Segment
X14208 N14208 N14209 Segment
X14209 N14209 N14210 Segment
X14210 N14210 N14211 Segment
X14211 N14211 N14212 Segment
X14212 N14212 N14213 Segment
X14213 N14213 N14214 Segment
X14214 N14214 N14215 Segment
X14215 N14215 N14216 Segment
X14216 N14216 N14217 Segment
X14217 N14217 N14218 Segment
X14218 N14218 N14219 Segment
X14219 N14219 N14220 Segment
X14220 N14220 N14221 Segment
X14221 N14221 N14222 Segment
X14222 N14222 N14223 Segment
X14223 N14223 N14224 Segment
X14224 N14224 N14225 Segment
X14225 N14225 N14226 Segment
X14226 N14226 N14227 Segment
X14227 N14227 N14228 Segment
X14228 N14228 N14229 Segment
X14229 N14229 N14230 Segment
X14230 N14230 N14231 Segment
X14231 N14231 N14232 Segment
X14232 N14232 N14233 Segment
X14233 N14233 N14234 Segment
X14234 N14234 N14235 Segment
X14235 N14235 N14236 Segment
X14236 N14236 N14237 Segment
X14237 N14237 N14238 Segment
X14238 N14238 N14239 Segment
X14239 N14239 N14240 Segment
X14240 N14240 N14241 Segment
X14241 N14241 N14242 Segment
X14242 N14242 N14243 Segment
X14243 N14243 N14244 Segment
X14244 N14244 N14245 Segment
X14245 N14245 N14246 Segment
X14246 N14246 N14247 Segment
X14247 N14247 N14248 Segment
X14248 N14248 N14249 Segment
X14249 N14249 N14250 Segment
X14250 N14250 N14251 Segment
X14251 N14251 N14252 Segment
X14252 N14252 N14253 Segment
X14253 N14253 N14254 Segment
X14254 N14254 N14255 Segment
X14255 N14255 N14256 Segment
X14256 N14256 N14257 Segment
X14257 N14257 N14258 Segment
X14258 N14258 N14259 Segment
X14259 N14259 N14260 Segment
X14260 N14260 N14261 Segment
X14261 N14261 N14262 Segment
X14262 N14262 N14263 Segment
X14263 N14263 N14264 Segment
X14264 N14264 N14265 Segment
X14265 N14265 N14266 Segment
X14266 N14266 N14267 Segment
X14267 N14267 N14268 Segment
X14268 N14268 N14269 Segment
X14269 N14269 N14270 Segment
X14270 N14270 N14271 Segment
X14271 N14271 N14272 Segment
X14272 N14272 N14273 Segment
X14273 N14273 N14274 Segment
X14274 N14274 N14275 Segment
X14275 N14275 N14276 Segment
X14276 N14276 N14277 Segment
X14277 N14277 N14278 Segment
X14278 N14278 N14279 Segment
X14279 N14279 N14280 Segment
X14280 N14280 N14281 Segment
X14281 N14281 N14282 Segment
X14282 N14282 N14283 Segment
X14283 N14283 N14284 Segment
X14284 N14284 N14285 Segment
X14285 N14285 N14286 Segment
X14286 N14286 N14287 Segment
X14287 N14287 N14288 Segment
X14288 N14288 N14289 Segment
X14289 N14289 N14290 Segment
X14290 N14290 N14291 Segment
X14291 N14291 N14292 Segment
X14292 N14292 N14293 Segment
X14293 N14293 N14294 Segment
X14294 N14294 N14295 Segment
X14295 N14295 N14296 Segment
X14296 N14296 N14297 Segment
X14297 N14297 N14298 Segment
X14298 N14298 N14299 Segment
X14299 N14299 N14300 Segment
X14300 N14300 N14301 Segment
X14301 N14301 N14302 Segment
X14302 N14302 N14303 Segment
X14303 N14303 N14304 Segment
X14304 N14304 N14305 Segment
X14305 N14305 N14306 Segment
X14306 N14306 N14307 Segment
X14307 N14307 N14308 Segment
X14308 N14308 N14309 Segment
X14309 N14309 N14310 Segment
X14310 N14310 N14311 Segment
X14311 N14311 N14312 Segment
X14312 N14312 N14313 Segment
X14313 N14313 N14314 Segment
X14314 N14314 N14315 Segment
X14315 N14315 N14316 Segment
X14316 N14316 N14317 Segment
X14317 N14317 N14318 Segment
X14318 N14318 N14319 Segment
X14319 N14319 N14320 Segment
X14320 N14320 N14321 Segment
X14321 N14321 N14322 Segment
X14322 N14322 N14323 Segment
X14323 N14323 N14324 Segment
X14324 N14324 N14325 Segment
X14325 N14325 N14326 Segment
X14326 N14326 N14327 Segment
X14327 N14327 N14328 Segment
X14328 N14328 N14329 Segment
X14329 N14329 N14330 Segment
X14330 N14330 N14331 Segment
X14331 N14331 N14332 Segment
X14332 N14332 N14333 Segment
X14333 N14333 N14334 Segment
X14334 N14334 N14335 Segment
X14335 N14335 N14336 Segment
X14336 N14336 N14337 Segment
X14337 N14337 N14338 Segment
X14338 N14338 N14339 Segment
X14339 N14339 N14340 Segment
X14340 N14340 N14341 Segment
X14341 N14341 N14342 Segment
X14342 N14342 N14343 Segment
X14343 N14343 N14344 Segment
X14344 N14344 N14345 Segment
X14345 N14345 N14346 Segment
X14346 N14346 N14347 Segment
X14347 N14347 N14348 Segment
X14348 N14348 N14349 Segment
X14349 N14349 N14350 Segment
X14350 N14350 N14351 Segment
X14351 N14351 N14352 Segment
X14352 N14352 N14353 Segment
X14353 N14353 N14354 Segment
X14354 N14354 N14355 Segment
X14355 N14355 N14356 Segment
X14356 N14356 N14357 Segment
X14357 N14357 N14358 Segment
X14358 N14358 N14359 Segment
X14359 N14359 N14360 Segment
X14360 N14360 N14361 Segment
X14361 N14361 N14362 Segment
X14362 N14362 N14363 Segment
X14363 N14363 N14364 Segment
X14364 N14364 N14365 Segment
X14365 N14365 N14366 Segment
X14366 N14366 N14367 Segment
X14367 N14367 N14368 Segment
X14368 N14368 N14369 Segment
X14369 N14369 N14370 Segment
X14370 N14370 N14371 Segment
X14371 N14371 N14372 Segment
X14372 N14372 N14373 Segment
X14373 N14373 N14374 Segment
X14374 N14374 N14375 Segment
X14375 N14375 N14376 Segment
X14376 N14376 N14377 Segment
X14377 N14377 N14378 Segment
X14378 N14378 N14379 Segment
X14379 N14379 N14380 Segment
X14380 N14380 N14381 Segment
X14381 N14381 N14382 Segment
X14382 N14382 N14383 Segment
X14383 N14383 N14384 Segment
X14384 N14384 N14385 Segment
X14385 N14385 N14386 Segment
X14386 N14386 N14387 Segment
X14387 N14387 N14388 Segment
X14388 N14388 N14389 Segment
X14389 N14389 N14390 Segment
X14390 N14390 N14391 Segment
X14391 N14391 N14392 Segment
X14392 N14392 N14393 Segment
X14393 N14393 N14394 Segment
X14394 N14394 N14395 Segment
X14395 N14395 N14396 Segment
X14396 N14396 N14397 Segment
X14397 N14397 N14398 Segment
X14398 N14398 N14399 Segment
X14399 N14399 N14400 Segment
X14400 N14400 N14401 Segment
X14401 N14401 N14402 Segment
X14402 N14402 N14403 Segment
X14403 N14403 N14404 Segment
X14404 N14404 N14405 Segment
X14405 N14405 N14406 Segment
X14406 N14406 N14407 Segment
X14407 N14407 N14408 Segment
X14408 N14408 N14409 Segment
X14409 N14409 N14410 Segment
X14410 N14410 N14411 Segment
X14411 N14411 N14412 Segment
X14412 N14412 N14413 Segment
X14413 N14413 N14414 Segment
X14414 N14414 N14415 Segment
X14415 N14415 N14416 Segment
X14416 N14416 N14417 Segment
X14417 N14417 N14418 Segment
X14418 N14418 N14419 Segment
X14419 N14419 N14420 Segment
X14420 N14420 N14421 Segment
X14421 N14421 N14422 Segment
X14422 N14422 N14423 Segment
X14423 N14423 N14424 Segment
X14424 N14424 N14425 Segment
X14425 N14425 N14426 Segment
X14426 N14426 N14427 Segment
X14427 N14427 N14428 Segment
X14428 N14428 N14429 Segment
X14429 N14429 N14430 Segment
X14430 N14430 N14431 Segment
X14431 N14431 N14432 Segment
X14432 N14432 N14433 Segment
X14433 N14433 N14434 Segment
X14434 N14434 N14435 Segment
X14435 N14435 N14436 Segment
X14436 N14436 N14437 Segment
X14437 N14437 N14438 Segment
X14438 N14438 N14439 Segment
X14439 N14439 N14440 Segment
X14440 N14440 N14441 Segment
X14441 N14441 N14442 Segment
X14442 N14442 N14443 Segment
X14443 N14443 N14444 Segment
X14444 N14444 N14445 Segment
X14445 N14445 N14446 Segment
X14446 N14446 N14447 Segment
X14447 N14447 N14448 Segment
X14448 N14448 N14449 Segment
X14449 N14449 N14450 Segment
X14450 N14450 N14451 Segment
X14451 N14451 N14452 Segment
X14452 N14452 N14453 Segment
X14453 N14453 N14454 Segment
X14454 N14454 N14455 Segment
X14455 N14455 N14456 Segment
X14456 N14456 N14457 Segment
X14457 N14457 N14458 Segment
X14458 N14458 N14459 Segment
X14459 N14459 N14460 Segment
X14460 N14460 N14461 Segment
X14461 N14461 N14462 Segment
X14462 N14462 N14463 Segment
X14463 N14463 N14464 Segment
X14464 N14464 N14465 Segment
X14465 N14465 N14466 Segment
X14466 N14466 N14467 Segment
X14467 N14467 N14468 Segment
X14468 N14468 N14469 Segment
X14469 N14469 N14470 Segment
X14470 N14470 N14471 Segment
X14471 N14471 N14472 Segment
X14472 N14472 N14473 Segment
X14473 N14473 N14474 Segment
X14474 N14474 N14475 Segment
X14475 N14475 N14476 Segment
X14476 N14476 N14477 Segment
X14477 N14477 N14478 Segment
X14478 N14478 N14479 Segment
X14479 N14479 N14480 Segment
X14480 N14480 N14481 Segment
X14481 N14481 N14482 Segment
X14482 N14482 N14483 Segment
X14483 N14483 N14484 Segment
X14484 N14484 N14485 Segment
X14485 N14485 N14486 Segment
X14486 N14486 N14487 Segment
X14487 N14487 N14488 Segment
X14488 N14488 N14489 Segment
X14489 N14489 N14490 Segment
X14490 N14490 N14491 Segment
X14491 N14491 N14492 Segment
X14492 N14492 N14493 Segment
X14493 N14493 N14494 Segment
X14494 N14494 N14495 Segment
X14495 N14495 N14496 Segment
X14496 N14496 N14497 Segment
X14497 N14497 N14498 Segment
X14498 N14498 N14499 Segment
X14499 N14499 N14500 Segment
X14500 N14500 N14501 Segment
X14501 N14501 N14502 Segment
X14502 N14502 N14503 Segment
X14503 N14503 N14504 Segment
X14504 N14504 N14505 Segment
X14505 N14505 N14506 Segment
X14506 N14506 N14507 Segment
X14507 N14507 N14508 Segment
X14508 N14508 N14509 Segment
X14509 N14509 N14510 Segment
X14510 N14510 N14511 Segment
X14511 N14511 N14512 Segment
X14512 N14512 N14513 Segment
X14513 N14513 N14514 Segment
X14514 N14514 N14515 Segment
X14515 N14515 N14516 Segment
X14516 N14516 N14517 Segment
X14517 N14517 N14518 Segment
X14518 N14518 N14519 Segment
X14519 N14519 N14520 Segment
X14520 N14520 N14521 Segment
X14521 N14521 N14522 Segment
X14522 N14522 N14523 Segment
X14523 N14523 N14524 Segment
X14524 N14524 N14525 Segment
X14525 N14525 N14526 Segment
X14526 N14526 N14527 Segment
X14527 N14527 N14528 Segment
X14528 N14528 N14529 Segment
X14529 N14529 N14530 Segment
X14530 N14530 N14531 Segment
X14531 N14531 N14532 Segment
X14532 N14532 N14533 Segment
X14533 N14533 N14534 Segment
X14534 N14534 N14535 Segment
X14535 N14535 N14536 Segment
X14536 N14536 N14537 Segment
X14537 N14537 N14538 Segment
X14538 N14538 N14539 Segment
X14539 N14539 N14540 Segment
X14540 N14540 N14541 Segment
X14541 N14541 N14542 Segment
X14542 N14542 N14543 Segment
X14543 N14543 N14544 Segment
X14544 N14544 N14545 Segment
X14545 N14545 N14546 Segment
X14546 N14546 N14547 Segment
X14547 N14547 N14548 Segment
X14548 N14548 N14549 Segment
X14549 N14549 N14550 Segment
X14550 N14550 N14551 Segment
X14551 N14551 N14552 Segment
X14552 N14552 N14553 Segment
X14553 N14553 N14554 Segment
X14554 N14554 N14555 Segment
X14555 N14555 N14556 Segment
X14556 N14556 N14557 Segment
X14557 N14557 N14558 Segment
X14558 N14558 N14559 Segment
X14559 N14559 N14560 Segment
X14560 N14560 N14561 Segment
X14561 N14561 N14562 Segment
X14562 N14562 N14563 Segment
X14563 N14563 N14564 Segment
X14564 N14564 N14565 Segment
X14565 N14565 N14566 Segment
X14566 N14566 N14567 Segment
X14567 N14567 N14568 Segment
X14568 N14568 N14569 Segment
X14569 N14569 N14570 Segment
X14570 N14570 N14571 Segment
X14571 N14571 N14572 Segment
X14572 N14572 N14573 Segment
X14573 N14573 N14574 Segment
X14574 N14574 N14575 Segment
X14575 N14575 N14576 Segment
X14576 N14576 N14577 Segment
X14577 N14577 N14578 Segment
X14578 N14578 N14579 Segment
X14579 N14579 N14580 Segment
X14580 N14580 N14581 Segment
X14581 N14581 N14582 Segment
X14582 N14582 N14583 Segment
X14583 N14583 N14584 Segment
X14584 N14584 N14585 Segment
X14585 N14585 N14586 Segment
X14586 N14586 N14587 Segment
X14587 N14587 N14588 Segment
X14588 N14588 N14589 Segment
X14589 N14589 N14590 Segment
X14590 N14590 N14591 Segment
X14591 N14591 N14592 Segment
X14592 N14592 N14593 Segment
X14593 N14593 N14594 Segment
X14594 N14594 N14595 Segment
X14595 N14595 N14596 Segment
X14596 N14596 N14597 Segment
X14597 N14597 N14598 Segment
X14598 N14598 N14599 Segment
X14599 N14599 N14600 Segment
X14600 N14600 N14601 Segment
X14601 N14601 N14602 Segment
X14602 N14602 N14603 Segment
X14603 N14603 N14604 Segment
X14604 N14604 N14605 Segment
X14605 N14605 N14606 Segment
X14606 N14606 N14607 Segment
X14607 N14607 N14608 Segment
X14608 N14608 N14609 Segment
X14609 N14609 N14610 Segment
X14610 N14610 N14611 Segment
X14611 N14611 N14612 Segment
X14612 N14612 N14613 Segment
X14613 N14613 N14614 Segment
X14614 N14614 N14615 Segment
X14615 N14615 N14616 Segment
X14616 N14616 N14617 Segment
X14617 N14617 N14618 Segment
X14618 N14618 N14619 Segment
X14619 N14619 N14620 Segment
X14620 N14620 N14621 Segment
X14621 N14621 N14622 Segment
X14622 N14622 N14623 Segment
X14623 N14623 N14624 Segment
X14624 N14624 N14625 Segment
X14625 N14625 N14626 Segment
X14626 N14626 N14627 Segment
X14627 N14627 N14628 Segment
X14628 N14628 N14629 Segment
X14629 N14629 N14630 Segment
X14630 N14630 N14631 Segment
X14631 N14631 N14632 Segment
X14632 N14632 N14633 Segment
X14633 N14633 N14634 Segment
X14634 N14634 N14635 Segment
X14635 N14635 N14636 Segment
X14636 N14636 N14637 Segment
X14637 N14637 N14638 Segment
X14638 N14638 N14639 Segment
X14639 N14639 N14640 Segment
X14640 N14640 N14641 Segment
X14641 N14641 N14642 Segment
X14642 N14642 N14643 Segment
X14643 N14643 N14644 Segment
X14644 N14644 N14645 Segment
X14645 N14645 N14646 Segment
X14646 N14646 N14647 Segment
X14647 N14647 N14648 Segment
X14648 N14648 N14649 Segment
X14649 N14649 N14650 Segment
X14650 N14650 N14651 Segment
X14651 N14651 N14652 Segment
X14652 N14652 N14653 Segment
X14653 N14653 N14654 Segment
X14654 N14654 N14655 Segment
X14655 N14655 N14656 Segment
X14656 N14656 N14657 Segment
X14657 N14657 N14658 Segment
X14658 N14658 N14659 Segment
X14659 N14659 N14660 Segment
X14660 N14660 N14661 Segment
X14661 N14661 N14662 Segment
X14662 N14662 N14663 Segment
X14663 N14663 N14664 Segment
X14664 N14664 N14665 Segment
X14665 N14665 N14666 Segment
X14666 N14666 N14667 Segment
X14667 N14667 N14668 Segment
X14668 N14668 N14669 Segment
X14669 N14669 N14670 Segment
X14670 N14670 N14671 Segment
X14671 N14671 N14672 Segment
X14672 N14672 N14673 Segment
X14673 N14673 N14674 Segment
X14674 N14674 N14675 Segment
X14675 N14675 N14676 Segment
X14676 N14676 N14677 Segment
X14677 N14677 N14678 Segment
X14678 N14678 N14679 Segment
X14679 N14679 N14680 Segment
X14680 N14680 N14681 Segment
X14681 N14681 N14682 Segment
X14682 N14682 N14683 Segment
X14683 N14683 N14684 Segment
X14684 N14684 N14685 Segment
X14685 N14685 N14686 Segment
X14686 N14686 N14687 Segment
X14687 N14687 N14688 Segment
X14688 N14688 N14689 Segment
X14689 N14689 N14690 Segment
X14690 N14690 N14691 Segment
X14691 N14691 N14692 Segment
X14692 N14692 N14693 Segment
X14693 N14693 N14694 Segment
X14694 N14694 N14695 Segment
X14695 N14695 N14696 Segment
X14696 N14696 N14697 Segment
X14697 N14697 N14698 Segment
X14698 N14698 N14699 Segment
X14699 N14699 N14700 Segment
X14700 N14700 N14701 Segment
X14701 N14701 N14702 Segment
X14702 N14702 N14703 Segment
X14703 N14703 N14704 Segment
X14704 N14704 N14705 Segment
X14705 N14705 N14706 Segment
X14706 N14706 N14707 Segment
X14707 N14707 N14708 Segment
X14708 N14708 N14709 Segment
X14709 N14709 N14710 Segment
X14710 N14710 N14711 Segment
X14711 N14711 N14712 Segment
X14712 N14712 N14713 Segment
X14713 N14713 N14714 Segment
X14714 N14714 N14715 Segment
X14715 N14715 N14716 Segment
X14716 N14716 N14717 Segment
X14717 N14717 N14718 Segment
X14718 N14718 N14719 Segment
X14719 N14719 N14720 Segment
X14720 N14720 N14721 Segment
X14721 N14721 N14722 Segment
X14722 N14722 N14723 Segment
X14723 N14723 N14724 Segment
X14724 N14724 N14725 Segment
X14725 N14725 N14726 Segment
X14726 N14726 N14727 Segment
X14727 N14727 N14728 Segment
X14728 N14728 N14729 Segment
X14729 N14729 N14730 Segment
X14730 N14730 N14731 Segment
X14731 N14731 N14732 Segment
X14732 N14732 N14733 Segment
X14733 N14733 N14734 Segment
X14734 N14734 N14735 Segment
X14735 N14735 N14736 Segment
X14736 N14736 N14737 Segment
X14737 N14737 N14738 Segment
X14738 N14738 N14739 Segment
X14739 N14739 N14740 Segment
X14740 N14740 N14741 Segment
X14741 N14741 N14742 Segment
X14742 N14742 N14743 Segment
X14743 N14743 N14744 Segment
X14744 N14744 N14745 Segment
X14745 N14745 N14746 Segment
X14746 N14746 N14747 Segment
X14747 N14747 N14748 Segment
X14748 N14748 N14749 Segment
X14749 N14749 N14750 Segment
X14750 N14750 N14751 Segment
X14751 N14751 N14752 Segment
X14752 N14752 N14753 Segment
X14753 N14753 N14754 Segment
X14754 N14754 N14755 Segment
X14755 N14755 N14756 Segment
X14756 N14756 N14757 Segment
X14757 N14757 N14758 Segment
X14758 N14758 N14759 Segment
X14759 N14759 N14760 Segment
X14760 N14760 N14761 Segment
X14761 N14761 N14762 Segment
X14762 N14762 N14763 Segment
X14763 N14763 N14764 Segment
X14764 N14764 N14765 Segment
X14765 N14765 N14766 Segment
X14766 N14766 N14767 Segment
X14767 N14767 N14768 Segment
X14768 N14768 N14769 Segment
X14769 N14769 N14770 Segment
X14770 N14770 N14771 Segment
X14771 N14771 N14772 Segment
X14772 N14772 N14773 Segment
X14773 N14773 N14774 Segment
X14774 N14774 N14775 Segment
X14775 N14775 N14776 Segment
X14776 N14776 N14777 Segment
X14777 N14777 N14778 Segment
X14778 N14778 N14779 Segment
X14779 N14779 N14780 Segment
X14780 N14780 N14781 Segment
X14781 N14781 N14782 Segment
X14782 N14782 N14783 Segment
X14783 N14783 N14784 Segment
X14784 N14784 N14785 Segment
X14785 N14785 N14786 Segment
X14786 N14786 N14787 Segment
X14787 N14787 N14788 Segment
X14788 N14788 N14789 Segment
X14789 N14789 N14790 Segment
X14790 N14790 N14791 Segment
X14791 N14791 N14792 Segment
X14792 N14792 N14793 Segment
X14793 N14793 N14794 Segment
X14794 N14794 N14795 Segment
X14795 N14795 N14796 Segment
X14796 N14796 N14797 Segment
X14797 N14797 N14798 Segment
X14798 N14798 N14799 Segment
X14799 N14799 N14800 Segment
X14800 N14800 N14801 Segment
X14801 N14801 N14802 Segment
X14802 N14802 N14803 Segment
X14803 N14803 N14804 Segment
X14804 N14804 N14805 Segment
X14805 N14805 N14806 Segment
X14806 N14806 N14807 Segment
X14807 N14807 N14808 Segment
X14808 N14808 N14809 Segment
X14809 N14809 N14810 Segment
X14810 N14810 N14811 Segment
X14811 N14811 N14812 Segment
X14812 N14812 N14813 Segment
X14813 N14813 N14814 Segment
X14814 N14814 N14815 Segment
X14815 N14815 N14816 Segment
X14816 N14816 N14817 Segment
X14817 N14817 N14818 Segment
X14818 N14818 N14819 Segment
X14819 N14819 N14820 Segment
X14820 N14820 N14821 Segment
X14821 N14821 N14822 Segment
X14822 N14822 N14823 Segment
X14823 N14823 N14824 Segment
X14824 N14824 N14825 Segment
X14825 N14825 N14826 Segment
X14826 N14826 N14827 Segment
X14827 N14827 N14828 Segment
X14828 N14828 N14829 Segment
X14829 N14829 N14830 Segment
X14830 N14830 N14831 Segment
X14831 N14831 N14832 Segment
X14832 N14832 N14833 Segment
X14833 N14833 N14834 Segment
X14834 N14834 N14835 Segment
X14835 N14835 N14836 Segment
X14836 N14836 N14837 Segment
X14837 N14837 N14838 Segment
X14838 N14838 N14839 Segment
X14839 N14839 N14840 Segment
X14840 N14840 N14841 Segment
X14841 N14841 N14842 Segment
X14842 N14842 N14843 Segment
X14843 N14843 N14844 Segment
X14844 N14844 N14845 Segment
X14845 N14845 N14846 Segment
X14846 N14846 N14847 Segment
X14847 N14847 N14848 Segment
X14848 N14848 N14849 Segment
X14849 N14849 N14850 Segment
X14850 N14850 N14851 Segment
X14851 N14851 N14852 Segment
X14852 N14852 N14853 Segment
X14853 N14853 N14854 Segment
X14854 N14854 N14855 Segment
X14855 N14855 N14856 Segment
X14856 N14856 N14857 Segment
X14857 N14857 N14858 Segment
X14858 N14858 N14859 Segment
X14859 N14859 N14860 Segment
X14860 N14860 N14861 Segment
X14861 N14861 N14862 Segment
X14862 N14862 N14863 Segment
X14863 N14863 N14864 Segment
X14864 N14864 N14865 Segment
X14865 N14865 N14866 Segment
X14866 N14866 N14867 Segment
X14867 N14867 N14868 Segment
X14868 N14868 N14869 Segment
X14869 N14869 N14870 Segment
X14870 N14870 N14871 Segment
X14871 N14871 N14872 Segment
X14872 N14872 N14873 Segment
X14873 N14873 N14874 Segment
X14874 N14874 N14875 Segment
X14875 N14875 N14876 Segment
X14876 N14876 N14877 Segment
X14877 N14877 N14878 Segment
X14878 N14878 N14879 Segment
X14879 N14879 N14880 Segment
X14880 N14880 N14881 Segment
X14881 N14881 N14882 Segment
X14882 N14882 N14883 Segment
X14883 N14883 N14884 Segment
X14884 N14884 N14885 Segment
X14885 N14885 N14886 Segment
X14886 N14886 N14887 Segment
X14887 N14887 N14888 Segment
X14888 N14888 N14889 Segment
X14889 N14889 N14890 Segment
X14890 N14890 N14891 Segment
X14891 N14891 N14892 Segment
X14892 N14892 N14893 Segment
X14893 N14893 N14894 Segment
X14894 N14894 N14895 Segment
X14895 N14895 N14896 Segment
X14896 N14896 N14897 Segment
X14897 N14897 N14898 Segment
X14898 N14898 N14899 Segment
X14899 N14899 N14900 Segment
X14900 N14900 N14901 Segment
X14901 N14901 N14902 Segment
X14902 N14902 N14903 Segment
X14903 N14903 N14904 Segment
X14904 N14904 N14905 Segment
X14905 N14905 N14906 Segment
X14906 N14906 N14907 Segment
X14907 N14907 N14908 Segment
X14908 N14908 N14909 Segment
X14909 N14909 N14910 Segment
X14910 N14910 N14911 Segment
X14911 N14911 N14912 Segment
X14912 N14912 N14913 Segment
X14913 N14913 N14914 Segment
X14914 N14914 N14915 Segment
X14915 N14915 N14916 Segment
X14916 N14916 N14917 Segment
X14917 N14917 N14918 Segment
X14918 N14918 N14919 Segment
X14919 N14919 N14920 Segment
X14920 N14920 N14921 Segment
X14921 N14921 N14922 Segment
X14922 N14922 N14923 Segment
X14923 N14923 N14924 Segment
X14924 N14924 N14925 Segment
X14925 N14925 N14926 Segment
X14926 N14926 N14927 Segment
X14927 N14927 N14928 Segment
X14928 N14928 N14929 Segment
X14929 N14929 N14930 Segment
X14930 N14930 N14931 Segment
X14931 N14931 N14932 Segment
X14932 N14932 N14933 Segment
X14933 N14933 N14934 Segment
X14934 N14934 N14935 Segment
X14935 N14935 N14936 Segment
X14936 N14936 N14937 Segment
X14937 N14937 N14938 Segment
X14938 N14938 N14939 Segment
X14939 N14939 N14940 Segment
X14940 N14940 N14941 Segment
X14941 N14941 N14942 Segment
X14942 N14942 N14943 Segment
X14943 N14943 N14944 Segment
X14944 N14944 N14945 Segment
X14945 N14945 N14946 Segment
X14946 N14946 N14947 Segment
X14947 N14947 N14948 Segment
X14948 N14948 N14949 Segment
X14949 N14949 N14950 Segment
X14950 N14950 N14951 Segment
X14951 N14951 N14952 Segment
X14952 N14952 N14953 Segment
X14953 N14953 N14954 Segment
X14954 N14954 N14955 Segment
X14955 N14955 N14956 Segment
X14956 N14956 N14957 Segment
X14957 N14957 N14958 Segment
X14958 N14958 N14959 Segment
X14959 N14959 N14960 Segment
X14960 N14960 N14961 Segment
X14961 N14961 N14962 Segment
X14962 N14962 N14963 Segment
X14963 N14963 N14964 Segment
X14964 N14964 N14965 Segment
X14965 N14965 N14966 Segment
X14966 N14966 N14967 Segment
X14967 N14967 N14968 Segment
X14968 N14968 N14969 Segment
X14969 N14969 N14970 Segment
X14970 N14970 N14971 Segment
X14971 N14971 N14972 Segment
X14972 N14972 N14973 Segment
X14973 N14973 N14974 Segment
X14974 N14974 N14975 Segment
X14975 N14975 N14976 Segment
X14976 N14976 N14977 Segment
X14977 N14977 N14978 Segment
X14978 N14978 N14979 Segment
X14979 N14979 N14980 Segment
X14980 N14980 N14981 Segment
X14981 N14981 N14982 Segment
X14982 N14982 N14983 Segment
X14983 N14983 N14984 Segment
X14984 N14984 N14985 Segment
X14985 N14985 N14986 Segment
X14986 N14986 N14987 Segment
X14987 N14987 N14988 Segment
X14988 N14988 N14989 Segment
X14989 N14989 N14990 Segment
X14990 N14990 N14991 Segment
X14991 N14991 N14992 Segment
X14992 N14992 N14993 Segment
X14993 N14993 N14994 Segment
X14994 N14994 N14995 Segment
X14995 N14995 N14996 Segment
X14996 N14996 N14997 Segment
X14997 N14997 N14998 Segment
X14998 N14998 N14999 Segment
X14999 N14999 N15000 Segment
X15000 N15000 N15001 Segment
X15001 N15001 N15002 Segment
X15002 N15002 N15003 Segment
X15003 N15003 N15004 Segment
X15004 N15004 N15005 Segment
X15005 N15005 N15006 Segment
X15006 N15006 N15007 Segment
X15007 N15007 N15008 Segment
X15008 N15008 N15009 Segment
X15009 N15009 N15010 Segment
X15010 N15010 N15011 Segment
X15011 N15011 N15012 Segment
X15012 N15012 N15013 Segment
X15013 N15013 N15014 Segment
X15014 N15014 N15015 Segment
X15015 N15015 N15016 Segment
X15016 N15016 N15017 Segment
X15017 N15017 N15018 Segment
X15018 N15018 N15019 Segment
X15019 N15019 N15020 Segment
X15020 N15020 N15021 Segment
X15021 N15021 N15022 Segment
X15022 N15022 N15023 Segment
X15023 N15023 N15024 Segment
X15024 N15024 N15025 Segment
X15025 N15025 N15026 Segment
X15026 N15026 N15027 Segment
X15027 N15027 N15028 Segment
X15028 N15028 N15029 Segment
X15029 N15029 N15030 Segment
X15030 N15030 N15031 Segment
X15031 N15031 N15032 Segment
X15032 N15032 N15033 Segment
X15033 N15033 N15034 Segment
X15034 N15034 N15035 Segment
X15035 N15035 N15036 Segment
X15036 N15036 N15037 Segment
X15037 N15037 N15038 Segment
X15038 N15038 N15039 Segment
X15039 N15039 N15040 Segment
X15040 N15040 N15041 Segment
X15041 N15041 N15042 Segment
X15042 N15042 N15043 Segment
X15043 N15043 N15044 Segment
X15044 N15044 N15045 Segment
X15045 N15045 N15046 Segment
X15046 N15046 N15047 Segment
X15047 N15047 N15048 Segment
X15048 N15048 N15049 Segment
X15049 N15049 N15050 Segment
X15050 N15050 N15051 Segment
X15051 N15051 N15052 Segment
X15052 N15052 N15053 Segment
X15053 N15053 N15054 Segment
X15054 N15054 N15055 Segment
X15055 N15055 N15056 Segment
X15056 N15056 N15057 Segment
X15057 N15057 N15058 Segment
X15058 N15058 N15059 Segment
X15059 N15059 N15060 Segment
X15060 N15060 N15061 Segment
X15061 N15061 N15062 Segment
X15062 N15062 N15063 Segment
X15063 N15063 N15064 Segment
X15064 N15064 N15065 Segment
X15065 N15065 N15066 Segment
X15066 N15066 N15067 Segment
X15067 N15067 N15068 Segment
X15068 N15068 N15069 Segment
X15069 N15069 N15070 Segment
X15070 N15070 N15071 Segment
X15071 N15071 N15072 Segment
X15072 N15072 N15073 Segment
X15073 N15073 N15074 Segment
X15074 N15074 N15075 Segment
X15075 N15075 N15076 Segment
X15076 N15076 N15077 Segment
X15077 N15077 N15078 Segment
X15078 N15078 N15079 Segment
X15079 N15079 N15080 Segment
X15080 N15080 N15081 Segment
X15081 N15081 N15082 Segment
X15082 N15082 N15083 Segment
X15083 N15083 N15084 Segment
X15084 N15084 N15085 Segment
X15085 N15085 N15086 Segment
X15086 N15086 N15087 Segment
X15087 N15087 N15088 Segment
X15088 N15088 N15089 Segment
X15089 N15089 N15090 Segment
X15090 N15090 N15091 Segment
X15091 N15091 N15092 Segment
X15092 N15092 N15093 Segment
X15093 N15093 N15094 Segment
X15094 N15094 N15095 Segment
X15095 N15095 N15096 Segment
X15096 N15096 N15097 Segment
X15097 N15097 N15098 Segment
X15098 N15098 N15099 Segment
X15099 N15099 N15100 Segment
X15100 N15100 N15101 Segment
X15101 N15101 N15102 Segment
X15102 N15102 N15103 Segment
X15103 N15103 N15104 Segment
X15104 N15104 N15105 Segment
X15105 N15105 N15106 Segment
X15106 N15106 N15107 Segment
X15107 N15107 N15108 Segment
X15108 N15108 N15109 Segment
X15109 N15109 N15110 Segment
X15110 N15110 N15111 Segment
X15111 N15111 N15112 Segment
X15112 N15112 N15113 Segment
X15113 N15113 N15114 Segment
X15114 N15114 N15115 Segment
X15115 N15115 N15116 Segment
X15116 N15116 N15117 Segment
X15117 N15117 N15118 Segment
X15118 N15118 N15119 Segment
X15119 N15119 N15120 Segment
X15120 N15120 N15121 Segment
X15121 N15121 N15122 Segment
X15122 N15122 N15123 Segment
X15123 N15123 N15124 Segment
X15124 N15124 N15125 Segment
X15125 N15125 N15126 Segment
X15126 N15126 N15127 Segment
X15127 N15127 N15128 Segment
X15128 N15128 N15129 Segment
X15129 N15129 N15130 Segment
X15130 N15130 N15131 Segment
X15131 N15131 N15132 Segment
X15132 N15132 N15133 Segment
X15133 N15133 N15134 Segment
X15134 N15134 N15135 Segment
X15135 N15135 N15136 Segment
X15136 N15136 N15137 Segment
X15137 N15137 N15138 Segment
X15138 N15138 N15139 Segment
X15139 N15139 N15140 Segment
X15140 N15140 N15141 Segment
X15141 N15141 N15142 Segment
X15142 N15142 N15143 Segment
X15143 N15143 N15144 Segment
X15144 N15144 N15145 Segment
X15145 N15145 N15146 Segment
X15146 N15146 N15147 Segment
X15147 N15147 N15148 Segment
X15148 N15148 N15149 Segment
X15149 N15149 N15150 Segment
X15150 N15150 N15151 Segment
X15151 N15151 N15152 Segment
X15152 N15152 N15153 Segment
X15153 N15153 N15154 Segment
X15154 N15154 N15155 Segment
X15155 N15155 N15156 Segment
X15156 N15156 N15157 Segment
X15157 N15157 N15158 Segment
X15158 N15158 N15159 Segment
X15159 N15159 N15160 Segment
X15160 N15160 N15161 Segment
X15161 N15161 N15162 Segment
X15162 N15162 N15163 Segment
X15163 N15163 N15164 Segment
X15164 N15164 N15165 Segment
X15165 N15165 N15166 Segment
X15166 N15166 N15167 Segment
X15167 N15167 N15168 Segment
X15168 N15168 N15169 Segment
X15169 N15169 N15170 Segment
X15170 N15170 N15171 Segment
X15171 N15171 N15172 Segment
X15172 N15172 N15173 Segment
X15173 N15173 N15174 Segment
X15174 N15174 N15175 Segment
X15175 N15175 N15176 Segment
X15176 N15176 N15177 Segment
X15177 N15177 N15178 Segment
X15178 N15178 N15179 Segment
X15179 N15179 N15180 Segment
X15180 N15180 N15181 Segment
X15181 N15181 N15182 Segment
X15182 N15182 N15183 Segment
X15183 N15183 N15184 Segment
X15184 N15184 N15185 Segment
X15185 N15185 N15186 Segment
X15186 N15186 N15187 Segment
X15187 N15187 N15188 Segment
X15188 N15188 N15189 Segment
X15189 N15189 N15190 Segment
X15190 N15190 N15191 Segment
X15191 N15191 N15192 Segment
X15192 N15192 N15193 Segment
X15193 N15193 N15194 Segment
X15194 N15194 N15195 Segment
X15195 N15195 N15196 Segment
X15196 N15196 N15197 Segment
X15197 N15197 N15198 Segment
X15198 N15198 N15199 Segment
X15199 N15199 N15200 Segment
X15200 N15200 N15201 Segment
X15201 N15201 N15202 Segment
X15202 N15202 N15203 Segment
X15203 N15203 N15204 Segment
X15204 N15204 N15205 Segment
X15205 N15205 N15206 Segment
X15206 N15206 N15207 Segment
X15207 N15207 N15208 Segment
X15208 N15208 N15209 Segment
X15209 N15209 N15210 Segment
X15210 N15210 N15211 Segment
X15211 N15211 N15212 Segment
X15212 N15212 N15213 Segment
X15213 N15213 N15214 Segment
X15214 N15214 N15215 Segment
X15215 N15215 N15216 Segment
X15216 N15216 N15217 Segment
X15217 N15217 N15218 Segment
X15218 N15218 N15219 Segment
X15219 N15219 N15220 Segment
X15220 N15220 N15221 Segment
X15221 N15221 N15222 Segment
X15222 N15222 N15223 Segment
X15223 N15223 N15224 Segment
X15224 N15224 N15225 Segment
X15225 N15225 N15226 Segment
X15226 N15226 N15227 Segment
X15227 N15227 N15228 Segment
X15228 N15228 N15229 Segment
X15229 N15229 N15230 Segment
X15230 N15230 N15231 Segment
X15231 N15231 N15232 Segment
X15232 N15232 N15233 Segment
X15233 N15233 N15234 Segment
X15234 N15234 N15235 Segment
X15235 N15235 N15236 Segment
X15236 N15236 N15237 Segment
X15237 N15237 N15238 Segment
X15238 N15238 N15239 Segment
X15239 N15239 N15240 Segment
X15240 N15240 N15241 Segment
X15241 N15241 N15242 Segment
X15242 N15242 N15243 Segment
X15243 N15243 N15244 Segment
X15244 N15244 N15245 Segment
X15245 N15245 N15246 Segment
X15246 N15246 N15247 Segment
X15247 N15247 N15248 Segment
X15248 N15248 N15249 Segment
X15249 N15249 N15250 Segment
X15250 N15250 N15251 Segment
X15251 N15251 N15252 Segment
X15252 N15252 N15253 Segment
X15253 N15253 N15254 Segment
X15254 N15254 N15255 Segment
X15255 N15255 N15256 Segment
X15256 N15256 N15257 Segment
X15257 N15257 N15258 Segment
X15258 N15258 N15259 Segment
X15259 N15259 N15260 Segment
X15260 N15260 N15261 Segment
X15261 N15261 N15262 Segment
X15262 N15262 N15263 Segment
X15263 N15263 N15264 Segment
X15264 N15264 N15265 Segment
X15265 N15265 N15266 Segment
X15266 N15266 N15267 Segment
X15267 N15267 N15268 Segment
X15268 N15268 N15269 Segment
X15269 N15269 N15270 Segment
X15270 N15270 N15271 Segment
X15271 N15271 N15272 Segment
X15272 N15272 N15273 Segment
X15273 N15273 N15274 Segment
X15274 N15274 N15275 Segment
X15275 N15275 N15276 Segment
X15276 N15276 N15277 Segment
X15277 N15277 N15278 Segment
X15278 N15278 N15279 Segment
X15279 N15279 N15280 Segment
X15280 N15280 N15281 Segment
X15281 N15281 N15282 Segment
X15282 N15282 N15283 Segment
X15283 N15283 N15284 Segment
X15284 N15284 N15285 Segment
X15285 N15285 N15286 Segment
X15286 N15286 N15287 Segment
X15287 N15287 N15288 Segment
X15288 N15288 N15289 Segment
X15289 N15289 N15290 Segment
X15290 N15290 N15291 Segment
X15291 N15291 N15292 Segment
X15292 N15292 N15293 Segment
X15293 N15293 N15294 Segment
X15294 N15294 N15295 Segment
X15295 N15295 N15296 Segment
X15296 N15296 N15297 Segment
X15297 N15297 N15298 Segment
X15298 N15298 N15299 Segment
X15299 N15299 N15300 Segment
X15300 N15300 N15301 Segment
X15301 N15301 N15302 Segment
X15302 N15302 N15303 Segment
X15303 N15303 N15304 Segment
X15304 N15304 N15305 Segment
X15305 N15305 N15306 Segment
X15306 N15306 N15307 Segment
X15307 N15307 N15308 Segment
X15308 N15308 N15309 Segment
X15309 N15309 N15310 Segment
X15310 N15310 N15311 Segment
X15311 N15311 N15312 Segment
X15312 N15312 N15313 Segment
X15313 N15313 N15314 Segment
X15314 N15314 N15315 Segment
X15315 N15315 N15316 Segment
X15316 N15316 N15317 Segment
X15317 N15317 N15318 Segment
X15318 N15318 N15319 Segment
X15319 N15319 N15320 Segment
X15320 N15320 N15321 Segment
X15321 N15321 N15322 Segment
X15322 N15322 N15323 Segment
X15323 N15323 N15324 Segment
X15324 N15324 N15325 Segment
X15325 N15325 N15326 Segment
X15326 N15326 N15327 Segment
X15327 N15327 N15328 Segment
X15328 N15328 N15329 Segment
X15329 N15329 N15330 Segment
X15330 N15330 N15331 Segment
X15331 N15331 N15332 Segment
X15332 N15332 N15333 Segment
X15333 N15333 N15334 Segment
X15334 N15334 N15335 Segment
X15335 N15335 N15336 Segment
X15336 N15336 N15337 Segment
X15337 N15337 N15338 Segment
X15338 N15338 N15339 Segment
X15339 N15339 N15340 Segment
X15340 N15340 N15341 Segment
X15341 N15341 N15342 Segment
X15342 N15342 N15343 Segment
X15343 N15343 N15344 Segment
X15344 N15344 N15345 Segment
X15345 N15345 N15346 Segment
X15346 N15346 N15347 Segment
X15347 N15347 N15348 Segment
X15348 N15348 N15349 Segment
X15349 N15349 N15350 Segment
X15350 N15350 N15351 Segment
X15351 N15351 N15352 Segment
X15352 N15352 N15353 Segment
X15353 N15353 N15354 Segment
X15354 N15354 N15355 Segment
X15355 N15355 N15356 Segment
X15356 N15356 N15357 Segment
X15357 N15357 N15358 Segment
X15358 N15358 N15359 Segment
X15359 N15359 N15360 Segment
X15360 N15360 N15361 Segment
X15361 N15361 N15362 Segment
X15362 N15362 N15363 Segment
X15363 N15363 N15364 Segment
X15364 N15364 N15365 Segment
X15365 N15365 N15366 Segment
X15366 N15366 N15367 Segment
X15367 N15367 N15368 Segment
X15368 N15368 N15369 Segment
X15369 N15369 N15370 Segment
X15370 N15370 N15371 Segment
X15371 N15371 N15372 Segment
X15372 N15372 N15373 Segment
X15373 N15373 N15374 Segment
X15374 N15374 N15375 Segment
X15375 N15375 N15376 Segment
X15376 N15376 N15377 Segment
X15377 N15377 N15378 Segment
X15378 N15378 N15379 Segment
X15379 N15379 N15380 Segment
X15380 N15380 N15381 Segment
X15381 N15381 N15382 Segment
X15382 N15382 N15383 Segment
X15383 N15383 N15384 Segment
X15384 N15384 N15385 Segment
X15385 N15385 N15386 Segment
X15386 N15386 N15387 Segment
X15387 N15387 N15388 Segment
X15388 N15388 N15389 Segment
X15389 N15389 N15390 Segment
X15390 N15390 N15391 Segment
X15391 N15391 N15392 Segment
X15392 N15392 N15393 Segment
X15393 N15393 N15394 Segment
X15394 N15394 N15395 Segment
X15395 N15395 N15396 Segment
X15396 N15396 N15397 Segment
X15397 N15397 N15398 Segment
X15398 N15398 N15399 Segment
X15399 N15399 N15400 Segment
X15400 N15400 N15401 Segment
X15401 N15401 N15402 Segment
X15402 N15402 N15403 Segment
X15403 N15403 N15404 Segment
X15404 N15404 N15405 Segment
X15405 N15405 N15406 Segment
X15406 N15406 N15407 Segment
X15407 N15407 N15408 Segment
X15408 N15408 N15409 Segment
X15409 N15409 N15410 Segment
X15410 N15410 N15411 Segment
X15411 N15411 N15412 Segment
X15412 N15412 N15413 Segment
X15413 N15413 N15414 Segment
X15414 N15414 N15415 Segment
X15415 N15415 N15416 Segment
X15416 N15416 N15417 Segment
X15417 N15417 N15418 Segment
X15418 N15418 N15419 Segment
X15419 N15419 N15420 Segment
X15420 N15420 N15421 Segment
X15421 N15421 N15422 Segment
X15422 N15422 N15423 Segment
X15423 N15423 N15424 Segment
X15424 N15424 N15425 Segment
X15425 N15425 N15426 Segment
X15426 N15426 N15427 Segment
X15427 N15427 N15428 Segment
X15428 N15428 N15429 Segment
X15429 N15429 N15430 Segment
X15430 N15430 N15431 Segment
X15431 N15431 N15432 Segment
X15432 N15432 N15433 Segment
X15433 N15433 N15434 Segment
X15434 N15434 N15435 Segment
X15435 N15435 N15436 Segment
X15436 N15436 N15437 Segment
X15437 N15437 N15438 Segment
X15438 N15438 N15439 Segment
X15439 N15439 N15440 Segment
X15440 N15440 N15441 Segment
X15441 N15441 N15442 Segment
X15442 N15442 N15443 Segment
X15443 N15443 N15444 Segment
X15444 N15444 N15445 Segment
X15445 N15445 N15446 Segment
X15446 N15446 N15447 Segment
X15447 N15447 N15448 Segment
X15448 N15448 N15449 Segment
X15449 N15449 N15450 Segment
X15450 N15450 N15451 Segment
X15451 N15451 N15452 Segment
X15452 N15452 N15453 Segment
X15453 N15453 N15454 Segment
X15454 N15454 N15455 Segment
X15455 N15455 N15456 Segment
X15456 N15456 N15457 Segment
X15457 N15457 N15458 Segment
X15458 N15458 N15459 Segment
X15459 N15459 N15460 Segment
X15460 N15460 N15461 Segment
X15461 N15461 N15462 Segment
X15462 N15462 N15463 Segment
X15463 N15463 N15464 Segment
X15464 N15464 N15465 Segment
X15465 N15465 N15466 Segment
X15466 N15466 N15467 Segment
X15467 N15467 N15468 Segment
X15468 N15468 N15469 Segment
X15469 N15469 N15470 Segment
X15470 N15470 N15471 Segment
X15471 N15471 N15472 Segment
X15472 N15472 N15473 Segment
X15473 N15473 N15474 Segment
X15474 N15474 N15475 Segment
X15475 N15475 N15476 Segment
X15476 N15476 N15477 Segment
X15477 N15477 N15478 Segment
X15478 N15478 N15479 Segment
X15479 N15479 N15480 Segment
X15480 N15480 N15481 Segment
X15481 N15481 N15482 Segment
X15482 N15482 N15483 Segment
X15483 N15483 N15484 Segment
X15484 N15484 N15485 Segment
X15485 N15485 N15486 Segment
X15486 N15486 N15487 Segment
X15487 N15487 N15488 Segment
X15488 N15488 N15489 Segment
X15489 N15489 N15490 Segment
X15490 N15490 N15491 Segment
X15491 N15491 N15492 Segment
X15492 N15492 N15493 Segment
X15493 N15493 N15494 Segment
X15494 N15494 N15495 Segment
X15495 N15495 N15496 Segment
X15496 N15496 N15497 Segment
X15497 N15497 N15498 Segment
X15498 N15498 N15499 Segment
X15499 N15499 N15500 Segment
X15500 N15500 N15501 Segment
X15501 N15501 N15502 Segment
X15502 N15502 N15503 Segment
X15503 N15503 N15504 Segment
X15504 N15504 N15505 Segment
X15505 N15505 N15506 Segment
X15506 N15506 N15507 Segment
X15507 N15507 N15508 Segment
X15508 N15508 N15509 Segment
X15509 N15509 N15510 Segment
X15510 N15510 N15511 Segment
X15511 N15511 N15512 Segment
X15512 N15512 N15513 Segment
X15513 N15513 N15514 Segment
X15514 N15514 N15515 Segment
X15515 N15515 N15516 Segment
X15516 N15516 N15517 Segment
X15517 N15517 N15518 Segment
X15518 N15518 N15519 Segment
X15519 N15519 N15520 Segment
X15520 N15520 N15521 Segment
X15521 N15521 N15522 Segment
X15522 N15522 N15523 Segment
X15523 N15523 N15524 Segment
X15524 N15524 N15525 Segment
X15525 N15525 N15526 Segment
X15526 N15526 N15527 Segment
X15527 N15527 N15528 Segment
X15528 N15528 N15529 Segment
X15529 N15529 N15530 Segment
X15530 N15530 N15531 Segment
X15531 N15531 N15532 Segment
X15532 N15532 N15533 Segment
X15533 N15533 N15534 Segment
X15534 N15534 N15535 Segment
X15535 N15535 N15536 Segment
X15536 N15536 N15537 Segment
X15537 N15537 N15538 Segment
X15538 N15538 N15539 Segment
X15539 N15539 N15540 Segment
X15540 N15540 N15541 Segment
X15541 N15541 N15542 Segment
X15542 N15542 N15543 Segment
X15543 N15543 N15544 Segment
X15544 N15544 N15545 Segment
X15545 N15545 N15546 Segment
X15546 N15546 N15547 Segment
X15547 N15547 N15548 Segment
X15548 N15548 N15549 Segment
X15549 N15549 N15550 Segment
X15550 N15550 N15551 Segment
X15551 N15551 N15552 Segment
X15552 N15552 N15553 Segment
X15553 N15553 N15554 Segment
X15554 N15554 N15555 Segment
X15555 N15555 N15556 Segment
X15556 N15556 N15557 Segment
X15557 N15557 N15558 Segment
X15558 N15558 N15559 Segment
X15559 N15559 N15560 Segment
X15560 N15560 N15561 Segment
X15561 N15561 N15562 Segment
X15562 N15562 N15563 Segment
X15563 N15563 N15564 Segment
X15564 N15564 N15565 Segment
X15565 N15565 N15566 Segment
X15566 N15566 N15567 Segment
X15567 N15567 N15568 Segment
X15568 N15568 N15569 Segment
X15569 N15569 N15570 Segment
X15570 N15570 N15571 Segment
X15571 N15571 N15572 Segment
X15572 N15572 N15573 Segment
X15573 N15573 N15574 Segment
X15574 N15574 N15575 Segment
X15575 N15575 N15576 Segment
X15576 N15576 N15577 Segment
X15577 N15577 N15578 Segment
X15578 N15578 N15579 Segment
X15579 N15579 N15580 Segment
X15580 N15580 N15581 Segment
X15581 N15581 N15582 Segment
X15582 N15582 N15583 Segment
X15583 N15583 N15584 Segment
X15584 N15584 N15585 Segment
X15585 N15585 N15586 Segment
X15586 N15586 N15587 Segment
X15587 N15587 N15588 Segment
X15588 N15588 N15589 Segment
X15589 N15589 N15590 Segment
X15590 N15590 N15591 Segment
X15591 N15591 N15592 Segment
X15592 N15592 N15593 Segment
X15593 N15593 N15594 Segment
X15594 N15594 N15595 Segment
X15595 N15595 N15596 Segment
X15596 N15596 N15597 Segment
X15597 N15597 N15598 Segment
X15598 N15598 N15599 Segment
X15599 N15599 N15600 Segment
X15600 N15600 N15601 Segment
X15601 N15601 N15602 Segment
X15602 N15602 N15603 Segment
X15603 N15603 N15604 Segment
X15604 N15604 N15605 Segment
X15605 N15605 N15606 Segment
X15606 N15606 N15607 Segment
X15607 N15607 N15608 Segment
X15608 N15608 N15609 Segment
X15609 N15609 N15610 Segment
X15610 N15610 N15611 Segment
X15611 N15611 N15612 Segment
X15612 N15612 N15613 Segment
X15613 N15613 N15614 Segment
X15614 N15614 N15615 Segment
X15615 N15615 N15616 Segment
X15616 N15616 N15617 Segment
X15617 N15617 N15618 Segment
X15618 N15618 N15619 Segment
X15619 N15619 N15620 Segment
X15620 N15620 N15621 Segment
X15621 N15621 N15622 Segment
X15622 N15622 N15623 Segment
X15623 N15623 N15624 Segment
X15624 N15624 N15625 Segment
X15625 N15625 N15626 Segment
X15626 N15626 N15627 Segment
X15627 N15627 N15628 Segment
X15628 N15628 N15629 Segment
X15629 N15629 N15630 Segment
X15630 N15630 N15631 Segment
X15631 N15631 N15632 Segment
X15632 N15632 N15633 Segment
X15633 N15633 N15634 Segment
X15634 N15634 N15635 Segment
X15635 N15635 N15636 Segment
X15636 N15636 N15637 Segment
X15637 N15637 N15638 Segment
X15638 N15638 N15639 Segment
X15639 N15639 N15640 Segment
X15640 N15640 N15641 Segment
X15641 N15641 N15642 Segment
X15642 N15642 N15643 Segment
X15643 N15643 N15644 Segment
X15644 N15644 N15645 Segment
X15645 N15645 N15646 Segment
X15646 N15646 N15647 Segment
X15647 N15647 N15648 Segment
X15648 N15648 N15649 Segment
X15649 N15649 N15650 Segment
X15650 N15650 N15651 Segment
X15651 N15651 N15652 Segment
X15652 N15652 N15653 Segment
X15653 N15653 N15654 Segment
X15654 N15654 N15655 Segment
X15655 N15655 N15656 Segment
X15656 N15656 N15657 Segment
X15657 N15657 N15658 Segment
X15658 N15658 N15659 Segment
X15659 N15659 N15660 Segment
X15660 N15660 N15661 Segment
X15661 N15661 N15662 Segment
X15662 N15662 N15663 Segment
X15663 N15663 N15664 Segment
X15664 N15664 N15665 Segment
X15665 N15665 N15666 Segment
X15666 N15666 N15667 Segment
X15667 N15667 N15668 Segment
X15668 N15668 N15669 Segment
X15669 N15669 N15670 Segment
X15670 N15670 N15671 Segment
X15671 N15671 N15672 Segment
X15672 N15672 N15673 Segment
X15673 N15673 N15674 Segment
X15674 N15674 N15675 Segment
X15675 N15675 N15676 Segment
X15676 N15676 N15677 Segment
X15677 N15677 N15678 Segment
X15678 N15678 N15679 Segment
X15679 N15679 N15680 Segment
X15680 N15680 N15681 Segment
X15681 N15681 N15682 Segment
X15682 N15682 N15683 Segment
X15683 N15683 N15684 Segment
X15684 N15684 N15685 Segment
X15685 N15685 N15686 Segment
X15686 N15686 N15687 Segment
X15687 N15687 N15688 Segment
X15688 N15688 N15689 Segment
X15689 N15689 N15690 Segment
X15690 N15690 N15691 Segment
X15691 N15691 N15692 Segment
X15692 N15692 N15693 Segment
X15693 N15693 N15694 Segment
X15694 N15694 N15695 Segment
X15695 N15695 N15696 Segment
X15696 N15696 N15697 Segment
X15697 N15697 N15698 Segment
X15698 N15698 N15699 Segment
X15699 N15699 N15700 Segment
X15700 N15700 N15701 Segment
X15701 N15701 N15702 Segment
X15702 N15702 N15703 Segment
X15703 N15703 N15704 Segment
X15704 N15704 N15705 Segment
X15705 N15705 N15706 Segment
X15706 N15706 N15707 Segment
X15707 N15707 N15708 Segment
X15708 N15708 N15709 Segment
X15709 N15709 N15710 Segment
X15710 N15710 N15711 Segment
X15711 N15711 N15712 Segment
X15712 N15712 N15713 Segment
X15713 N15713 N15714 Segment
X15714 N15714 N15715 Segment
X15715 N15715 N15716 Segment
X15716 N15716 N15717 Segment
X15717 N15717 N15718 Segment
X15718 N15718 N15719 Segment
X15719 N15719 N15720 Segment
X15720 N15720 N15721 Segment
X15721 N15721 N15722 Segment
X15722 N15722 N15723 Segment
X15723 N15723 N15724 Segment
X15724 N15724 N15725 Segment
X15725 N15725 N15726 Segment
X15726 N15726 N15727 Segment
X15727 N15727 N15728 Segment
X15728 N15728 N15729 Segment
X15729 N15729 N15730 Segment
X15730 N15730 N15731 Segment
X15731 N15731 N15732 Segment
X15732 N15732 N15733 Segment
X15733 N15733 N15734 Segment
X15734 N15734 N15735 Segment
X15735 N15735 N15736 Segment
X15736 N15736 N15737 Segment
X15737 N15737 N15738 Segment
X15738 N15738 N15739 Segment
X15739 N15739 N15740 Segment
X15740 N15740 N15741 Segment
X15741 N15741 N15742 Segment
X15742 N15742 N15743 Segment
X15743 N15743 N15744 Segment
X15744 N15744 N15745 Segment
X15745 N15745 N15746 Segment
X15746 N15746 N15747 Segment
X15747 N15747 N15748 Segment
X15748 N15748 N15749 Segment
X15749 N15749 N15750 Segment
X15750 N15750 N15751 Segment
X15751 N15751 N15752 Segment
X15752 N15752 N15753 Segment
X15753 N15753 N15754 Segment
X15754 N15754 N15755 Segment
X15755 N15755 N15756 Segment
X15756 N15756 N15757 Segment
X15757 N15757 N15758 Segment
X15758 N15758 N15759 Segment
X15759 N15759 N15760 Segment
X15760 N15760 N15761 Segment
X15761 N15761 N15762 Segment
X15762 N15762 N15763 Segment
X15763 N15763 N15764 Segment
X15764 N15764 N15765 Segment
X15765 N15765 N15766 Segment
X15766 N15766 N15767 Segment
X15767 N15767 N15768 Segment
X15768 N15768 N15769 Segment
X15769 N15769 N15770 Segment
X15770 N15770 N15771 Segment
X15771 N15771 N15772 Segment
X15772 N15772 N15773 Segment
X15773 N15773 N15774 Segment
X15774 N15774 N15775 Segment
X15775 N15775 N15776 Segment
X15776 N15776 N15777 Segment
X15777 N15777 N15778 Segment
X15778 N15778 N15779 Segment
X15779 N15779 N15780 Segment
X15780 N15780 N15781 Segment
X15781 N15781 N15782 Segment
X15782 N15782 N15783 Segment
X15783 N15783 N15784 Segment
X15784 N15784 N15785 Segment
X15785 N15785 N15786 Segment
X15786 N15786 N15787 Segment
X15787 N15787 N15788 Segment
X15788 N15788 N15789 Segment
X15789 N15789 N15790 Segment
X15790 N15790 N15791 Segment
X15791 N15791 N15792 Segment
X15792 N15792 N15793 Segment
X15793 N15793 N15794 Segment
X15794 N15794 N15795 Segment
X15795 N15795 N15796 Segment
X15796 N15796 N15797 Segment
X15797 N15797 N15798 Segment
X15798 N15798 N15799 Segment
X15799 N15799 N15800 Segment
X15800 N15800 N15801 Segment
X15801 N15801 N15802 Segment
X15802 N15802 N15803 Segment
X15803 N15803 N15804 Segment
X15804 N15804 N15805 Segment
X15805 N15805 N15806 Segment
X15806 N15806 N15807 Segment
X15807 N15807 N15808 Segment
X15808 N15808 N15809 Segment
X15809 N15809 N15810 Segment
X15810 N15810 N15811 Segment
X15811 N15811 N15812 Segment
X15812 N15812 N15813 Segment
X15813 N15813 N15814 Segment
X15814 N15814 N15815 Segment
X15815 N15815 N15816 Segment
X15816 N15816 N15817 Segment
X15817 N15817 N15818 Segment
X15818 N15818 N15819 Segment
X15819 N15819 N15820 Segment
X15820 N15820 N15821 Segment
X15821 N15821 N15822 Segment
X15822 N15822 N15823 Segment
X15823 N15823 N15824 Segment
X15824 N15824 N15825 Segment
X15825 N15825 N15826 Segment
X15826 N15826 N15827 Segment
X15827 N15827 N15828 Segment
X15828 N15828 N15829 Segment
X15829 N15829 N15830 Segment
X15830 N15830 N15831 Segment
X15831 N15831 N15832 Segment
X15832 N15832 N15833 Segment
X15833 N15833 N15834 Segment
X15834 N15834 N15835 Segment
X15835 N15835 N15836 Segment
X15836 N15836 N15837 Segment
X15837 N15837 N15838 Segment
X15838 N15838 N15839 Segment
X15839 N15839 N15840 Segment
X15840 N15840 N15841 Segment
X15841 N15841 N15842 Segment
X15842 N15842 N15843 Segment
X15843 N15843 N15844 Segment
X15844 N15844 N15845 Segment
X15845 N15845 N15846 Segment
X15846 N15846 N15847 Segment
X15847 N15847 N15848 Segment
X15848 N15848 N15849 Segment
X15849 N15849 N15850 Segment
X15850 N15850 N15851 Segment
X15851 N15851 N15852 Segment
X15852 N15852 N15853 Segment
X15853 N15853 N15854 Segment
X15854 N15854 N15855 Segment
X15855 N15855 N15856 Segment
X15856 N15856 N15857 Segment
X15857 N15857 N15858 Segment
X15858 N15858 N15859 Segment
X15859 N15859 N15860 Segment
X15860 N15860 N15861 Segment
X15861 N15861 N15862 Segment
X15862 N15862 N15863 Segment
X15863 N15863 N15864 Segment
X15864 N15864 N15865 Segment
X15865 N15865 N15866 Segment
X15866 N15866 N15867 Segment
X15867 N15867 N15868 Segment
X15868 N15868 N15869 Segment
X15869 N15869 N15870 Segment
X15870 N15870 N15871 Segment
X15871 N15871 N15872 Segment
X15872 N15872 N15873 Segment
X15873 N15873 N15874 Segment
X15874 N15874 N15875 Segment
X15875 N15875 N15876 Segment
X15876 N15876 N15877 Segment
X15877 N15877 N15878 Segment
X15878 N15878 N15879 Segment
X15879 N15879 N15880 Segment
X15880 N15880 N15881 Segment
X15881 N15881 N15882 Segment
X15882 N15882 N15883 Segment
X15883 N15883 N15884 Segment
X15884 N15884 N15885 Segment
X15885 N15885 N15886 Segment
X15886 N15886 N15887 Segment
X15887 N15887 N15888 Segment
X15888 N15888 N15889 Segment
X15889 N15889 N15890 Segment
X15890 N15890 N15891 Segment
X15891 N15891 N15892 Segment
X15892 N15892 N15893 Segment
X15893 N15893 N15894 Segment
X15894 N15894 N15895 Segment
X15895 N15895 N15896 Segment
X15896 N15896 N15897 Segment
X15897 N15897 N15898 Segment
X15898 N15898 N15899 Segment
X15899 N15899 N15900 Segment
X15900 N15900 N15901 Segment
X15901 N15901 N15902 Segment
X15902 N15902 N15903 Segment
X15903 N15903 N15904 Segment
X15904 N15904 N15905 Segment
X15905 N15905 N15906 Segment
X15906 N15906 N15907 Segment
X15907 N15907 N15908 Segment
X15908 N15908 N15909 Segment
X15909 N15909 N15910 Segment
X15910 N15910 N15911 Segment
X15911 N15911 N15912 Segment
X15912 N15912 N15913 Segment
X15913 N15913 N15914 Segment
X15914 N15914 N15915 Segment
X15915 N15915 N15916 Segment
X15916 N15916 N15917 Segment
X15917 N15917 N15918 Segment
X15918 N15918 N15919 Segment
X15919 N15919 N15920 Segment
X15920 N15920 N15921 Segment
X15921 N15921 N15922 Segment
X15922 N15922 N15923 Segment
X15923 N15923 N15924 Segment
X15924 N15924 N15925 Segment
X15925 N15925 N15926 Segment
X15926 N15926 N15927 Segment
X15927 N15927 N15928 Segment
X15928 N15928 N15929 Segment
X15929 N15929 N15930 Segment
X15930 N15930 N15931 Segment
X15931 N15931 N15932 Segment
X15932 N15932 N15933 Segment
X15933 N15933 N15934 Segment
X15934 N15934 N15935 Segment
X15935 N15935 N15936 Segment
X15936 N15936 N15937 Segment
X15937 N15937 N15938 Segment
X15938 N15938 N15939 Segment
X15939 N15939 N15940 Segment
X15940 N15940 N15941 Segment
X15941 N15941 N15942 Segment
X15942 N15942 N15943 Segment
X15943 N15943 N15944 Segment
X15944 N15944 N15945 Segment
X15945 N15945 N15946 Segment
X15946 N15946 N15947 Segment
X15947 N15947 N15948 Segment
X15948 N15948 N15949 Segment
X15949 N15949 N15950 Segment
X15950 N15950 N15951 Segment
X15951 N15951 N15952 Segment
X15952 N15952 N15953 Segment
X15953 N15953 N15954 Segment
X15954 N15954 N15955 Segment
X15955 N15955 N15956 Segment
X15956 N15956 N15957 Segment
X15957 N15957 N15958 Segment
X15958 N15958 N15959 Segment
X15959 N15959 N15960 Segment
X15960 N15960 N15961 Segment
X15961 N15961 N15962 Segment
X15962 N15962 N15963 Segment
X15963 N15963 N15964 Segment
X15964 N15964 N15965 Segment
X15965 N15965 N15966 Segment
X15966 N15966 N15967 Segment
X15967 N15967 N15968 Segment
X15968 N15968 N15969 Segment
X15969 N15969 N15970 Segment
X15970 N15970 N15971 Segment
X15971 N15971 N15972 Segment
X15972 N15972 N15973 Segment
X15973 N15973 N15974 Segment
X15974 N15974 N15975 Segment
X15975 N15975 N15976 Segment
X15976 N15976 N15977 Segment
X15977 N15977 N15978 Segment
X15978 N15978 N15979 Segment
X15979 N15979 N15980 Segment
X15980 N15980 N15981 Segment
X15981 N15981 N15982 Segment
X15982 N15982 N15983 Segment
X15983 N15983 N15984 Segment
X15984 N15984 N15985 Segment
X15985 N15985 N15986 Segment
X15986 N15986 N15987 Segment
X15987 N15987 N15988 Segment
X15988 N15988 N15989 Segment
X15989 N15989 N15990 Segment
X15990 N15990 N15991 Segment
X15991 N15991 N15992 Segment
X15992 N15992 N15993 Segment
X15993 N15993 N15994 Segment
X15994 N15994 N15995 Segment
X15995 N15995 N15996 Segment
X15996 N15996 N15997 Segment
X15997 N15997 N15998 Segment
X15998 N15998 N15999 Segment
X15999 N15999 N16000 Segment
X16000 N16000 N16001 Segment
X16001 N16001 N16002 Segment
X16002 N16002 N16003 Segment
X16003 N16003 N16004 Segment
X16004 N16004 N16005 Segment
X16005 N16005 N16006 Segment
X16006 N16006 N16007 Segment
X16007 N16007 N16008 Segment
X16008 N16008 N16009 Segment
X16009 N16009 N16010 Segment
X16010 N16010 N16011 Segment
X16011 N16011 N16012 Segment
X16012 N16012 N16013 Segment
X16013 N16013 N16014 Segment
X16014 N16014 N16015 Segment
X16015 N16015 N16016 Segment
X16016 N16016 N16017 Segment
X16017 N16017 N16018 Segment
X16018 N16018 N16019 Segment
X16019 N16019 N16020 Segment
X16020 N16020 N16021 Segment
X16021 N16021 N16022 Segment
X16022 N16022 N16023 Segment
X16023 N16023 N16024 Segment
X16024 N16024 N16025 Segment
X16025 N16025 N16026 Segment
X16026 N16026 N16027 Segment
X16027 N16027 N16028 Segment
X16028 N16028 N16029 Segment
X16029 N16029 N16030 Segment
X16030 N16030 N16031 Segment
X16031 N16031 N16032 Segment
X16032 N16032 N16033 Segment
X16033 N16033 N16034 Segment
X16034 N16034 N16035 Segment
X16035 N16035 N16036 Segment
X16036 N16036 N16037 Segment
X16037 N16037 N16038 Segment
X16038 N16038 N16039 Segment
X16039 N16039 N16040 Segment
X16040 N16040 N16041 Segment
X16041 N16041 N16042 Segment
X16042 N16042 N16043 Segment
X16043 N16043 N16044 Segment
X16044 N16044 N16045 Segment
X16045 N16045 N16046 Segment
X16046 N16046 N16047 Segment
X16047 N16047 N16048 Segment
X16048 N16048 N16049 Segment
X16049 N16049 N16050 Segment
X16050 N16050 N16051 Segment
X16051 N16051 N16052 Segment
X16052 N16052 N16053 Segment
X16053 N16053 N16054 Segment
X16054 N16054 N16055 Segment
X16055 N16055 N16056 Segment
X16056 N16056 N16057 Segment
X16057 N16057 N16058 Segment
X16058 N16058 N16059 Segment
X16059 N16059 N16060 Segment
X16060 N16060 N16061 Segment
X16061 N16061 N16062 Segment
X16062 N16062 N16063 Segment
X16063 N16063 N16064 Segment
X16064 N16064 N16065 Segment
X16065 N16065 N16066 Segment
X16066 N16066 N16067 Segment
X16067 N16067 N16068 Segment
X16068 N16068 N16069 Segment
X16069 N16069 N16070 Segment
X16070 N16070 N16071 Segment
X16071 N16071 N16072 Segment
X16072 N16072 N16073 Segment
X16073 N16073 N16074 Segment
X16074 N16074 N16075 Segment
X16075 N16075 N16076 Segment
X16076 N16076 N16077 Segment
X16077 N16077 N16078 Segment
X16078 N16078 N16079 Segment
X16079 N16079 N16080 Segment
X16080 N16080 N16081 Segment
X16081 N16081 N16082 Segment
X16082 N16082 N16083 Segment
X16083 N16083 N16084 Segment
X16084 N16084 N16085 Segment
X16085 N16085 N16086 Segment
X16086 N16086 N16087 Segment
X16087 N16087 N16088 Segment
X16088 N16088 N16089 Segment
X16089 N16089 N16090 Segment
X16090 N16090 N16091 Segment
X16091 N16091 N16092 Segment
X16092 N16092 N16093 Segment
X16093 N16093 N16094 Segment
X16094 N16094 N16095 Segment
X16095 N16095 N16096 Segment
X16096 N16096 N16097 Segment
X16097 N16097 N16098 Segment
X16098 N16098 N16099 Segment
X16099 N16099 N16100 Segment
X16100 N16100 N16101 Segment
X16101 N16101 N16102 Segment
X16102 N16102 N16103 Segment
X16103 N16103 N16104 Segment
X16104 N16104 N16105 Segment
X16105 N16105 N16106 Segment
X16106 N16106 N16107 Segment
X16107 N16107 N16108 Segment
X16108 N16108 N16109 Segment
X16109 N16109 N16110 Segment
X16110 N16110 N16111 Segment
X16111 N16111 N16112 Segment
X16112 N16112 N16113 Segment
X16113 N16113 N16114 Segment
X16114 N16114 N16115 Segment
X16115 N16115 N16116 Segment
X16116 N16116 N16117 Segment
X16117 N16117 N16118 Segment
X16118 N16118 N16119 Segment
X16119 N16119 N16120 Segment
X16120 N16120 N16121 Segment
X16121 N16121 N16122 Segment
X16122 N16122 N16123 Segment
X16123 N16123 N16124 Segment
X16124 N16124 N16125 Segment
X16125 N16125 N16126 Segment
X16126 N16126 N16127 Segment
X16127 N16127 N16128 Segment
X16128 N16128 N16129 Segment
X16129 N16129 N16130 Segment
X16130 N16130 N16131 Segment
X16131 N16131 N16132 Segment
X16132 N16132 N16133 Segment
X16133 N16133 N16134 Segment
X16134 N16134 N16135 Segment
X16135 N16135 N16136 Segment
X16136 N16136 N16137 Segment
X16137 N16137 N16138 Segment
X16138 N16138 N16139 Segment
X16139 N16139 N16140 Segment
X16140 N16140 N16141 Segment
X16141 N16141 N16142 Segment
X16142 N16142 N16143 Segment
X16143 N16143 N16144 Segment
X16144 N16144 N16145 Segment
X16145 N16145 N16146 Segment
X16146 N16146 N16147 Segment
X16147 N16147 N16148 Segment
X16148 N16148 N16149 Segment
X16149 N16149 N16150 Segment
X16150 N16150 N16151 Segment
X16151 N16151 N16152 Segment
X16152 N16152 N16153 Segment
X16153 N16153 N16154 Segment
X16154 N16154 N16155 Segment
X16155 N16155 N16156 Segment
X16156 N16156 N16157 Segment
X16157 N16157 N16158 Segment
X16158 N16158 N16159 Segment
X16159 N16159 N16160 Segment
X16160 N16160 N16161 Segment
X16161 N16161 N16162 Segment
X16162 N16162 N16163 Segment
X16163 N16163 N16164 Segment
X16164 N16164 N16165 Segment
X16165 N16165 N16166 Segment
X16166 N16166 N16167 Segment
X16167 N16167 N16168 Segment
X16168 N16168 N16169 Segment
X16169 N16169 N16170 Segment
X16170 N16170 N16171 Segment
X16171 N16171 N16172 Segment
X16172 N16172 N16173 Segment
X16173 N16173 N16174 Segment
X16174 N16174 N16175 Segment
X16175 N16175 N16176 Segment
X16176 N16176 N16177 Segment
X16177 N16177 N16178 Segment
X16178 N16178 N16179 Segment
X16179 N16179 N16180 Segment
X16180 N16180 N16181 Segment
X16181 N16181 N16182 Segment
X16182 N16182 N16183 Segment
X16183 N16183 N16184 Segment
X16184 N16184 N16185 Segment
X16185 N16185 N16186 Segment
X16186 N16186 N16187 Segment
X16187 N16187 N16188 Segment
X16188 N16188 N16189 Segment
X16189 N16189 N16190 Segment
X16190 N16190 N16191 Segment
X16191 N16191 N16192 Segment
X16192 N16192 N16193 Segment
X16193 N16193 N16194 Segment
X16194 N16194 N16195 Segment
X16195 N16195 N16196 Segment
X16196 N16196 N16197 Segment
X16197 N16197 N16198 Segment
X16198 N16198 N16199 Segment
X16199 N16199 N16200 Segment
X16200 N16200 N16201 Segment
X16201 N16201 N16202 Segment
X16202 N16202 N16203 Segment
X16203 N16203 N16204 Segment
X16204 N16204 N16205 Segment
X16205 N16205 N16206 Segment
X16206 N16206 N16207 Segment
X16207 N16207 N16208 Segment
X16208 N16208 N16209 Segment
X16209 N16209 N16210 Segment
X16210 N16210 N16211 Segment
X16211 N16211 N16212 Segment
X16212 N16212 N16213 Segment
X16213 N16213 N16214 Segment
X16214 N16214 N16215 Segment
X16215 N16215 N16216 Segment
X16216 N16216 N16217 Segment
X16217 N16217 N16218 Segment
X16218 N16218 N16219 Segment
X16219 N16219 N16220 Segment
X16220 N16220 N16221 Segment
X16221 N16221 N16222 Segment
X16222 N16222 N16223 Segment
X16223 N16223 N16224 Segment
X16224 N16224 N16225 Segment
X16225 N16225 N16226 Segment
X16226 N16226 N16227 Segment
X16227 N16227 N16228 Segment
X16228 N16228 N16229 Segment
X16229 N16229 N16230 Segment
X16230 N16230 N16231 Segment
X16231 N16231 N16232 Segment
X16232 N16232 N16233 Segment
X16233 N16233 N16234 Segment
X16234 N16234 N16235 Segment
X16235 N16235 N16236 Segment
X16236 N16236 N16237 Segment
X16237 N16237 N16238 Segment
X16238 N16238 N16239 Segment
X16239 N16239 N16240 Segment
X16240 N16240 N16241 Segment
X16241 N16241 N16242 Segment
X16242 N16242 N16243 Segment
X16243 N16243 N16244 Segment
X16244 N16244 N16245 Segment
X16245 N16245 N16246 Segment
X16246 N16246 N16247 Segment
X16247 N16247 N16248 Segment
X16248 N16248 N16249 Segment
X16249 N16249 N16250 Segment
X16250 N16250 N16251 Segment
X16251 N16251 N16252 Segment
X16252 N16252 N16253 Segment
X16253 N16253 N16254 Segment
X16254 N16254 N16255 Segment
X16255 N16255 N16256 Segment
X16256 N16256 N16257 Segment
X16257 N16257 N16258 Segment
X16258 N16258 N16259 Segment
X16259 N16259 N16260 Segment
X16260 N16260 N16261 Segment
X16261 N16261 N16262 Segment
X16262 N16262 N16263 Segment
X16263 N16263 N16264 Segment
X16264 N16264 N16265 Segment
X16265 N16265 N16266 Segment
X16266 N16266 N16267 Segment
X16267 N16267 N16268 Segment
X16268 N16268 N16269 Segment
X16269 N16269 N16270 Segment
X16270 N16270 N16271 Segment
X16271 N16271 N16272 Segment
X16272 N16272 N16273 Segment
X16273 N16273 N16274 Segment
X16274 N16274 N16275 Segment
X16275 N16275 N16276 Segment
X16276 N16276 N16277 Segment
X16277 N16277 N16278 Segment
X16278 N16278 N16279 Segment
X16279 N16279 N16280 Segment
X16280 N16280 N16281 Segment
X16281 N16281 N16282 Segment
X16282 N16282 N16283 Segment
X16283 N16283 N16284 Segment
X16284 N16284 N16285 Segment
X16285 N16285 N16286 Segment
X16286 N16286 N16287 Segment
X16287 N16287 N16288 Segment
X16288 N16288 N16289 Segment
X16289 N16289 N16290 Segment
X16290 N16290 N16291 Segment
X16291 N16291 N16292 Segment
X16292 N16292 N16293 Segment
X16293 N16293 N16294 Segment
X16294 N16294 N16295 Segment
X16295 N16295 N16296 Segment
X16296 N16296 N16297 Segment
X16297 N16297 N16298 Segment
X16298 N16298 N16299 Segment
X16299 N16299 N16300 Segment
X16300 N16300 N16301 Segment
X16301 N16301 N16302 Segment
X16302 N16302 N16303 Segment
X16303 N16303 N16304 Segment
X16304 N16304 N16305 Segment
X16305 N16305 N16306 Segment
X16306 N16306 N16307 Segment
X16307 N16307 N16308 Segment
X16308 N16308 N16309 Segment
X16309 N16309 N16310 Segment
X16310 N16310 N16311 Segment
X16311 N16311 N16312 Segment
X16312 N16312 N16313 Segment
X16313 N16313 N16314 Segment
X16314 N16314 N16315 Segment
X16315 N16315 N16316 Segment
X16316 N16316 N16317 Segment
X16317 N16317 N16318 Segment
X16318 N16318 N16319 Segment
X16319 N16319 N16320 Segment
X16320 N16320 N16321 Segment
X16321 N16321 N16322 Segment
X16322 N16322 N16323 Segment
X16323 N16323 N16324 Segment
X16324 N16324 N16325 Segment
X16325 N16325 N16326 Segment
X16326 N16326 N16327 Segment
X16327 N16327 N16328 Segment
X16328 N16328 N16329 Segment
X16329 N16329 N16330 Segment
X16330 N16330 N16331 Segment
X16331 N16331 N16332 Segment
X16332 N16332 N16333 Segment
X16333 N16333 N16334 Segment
X16334 N16334 N16335 Segment
X16335 N16335 N16336 Segment
X16336 N16336 N16337 Segment
X16337 N16337 N16338 Segment
X16338 N16338 N16339 Segment
X16339 N16339 N16340 Segment
X16340 N16340 N16341 Segment
X16341 N16341 N16342 Segment
X16342 N16342 N16343 Segment
X16343 N16343 N16344 Segment
X16344 N16344 N16345 Segment
X16345 N16345 N16346 Segment
X16346 N16346 N16347 Segment
X16347 N16347 N16348 Segment
X16348 N16348 N16349 Segment
X16349 N16349 N16350 Segment
X16350 N16350 N16351 Segment
X16351 N16351 N16352 Segment
X16352 N16352 N16353 Segment
X16353 N16353 N16354 Segment
X16354 N16354 N16355 Segment
X16355 N16355 N16356 Segment
X16356 N16356 N16357 Segment
X16357 N16357 N16358 Segment
X16358 N16358 N16359 Segment
X16359 N16359 N16360 Segment
X16360 N16360 N16361 Segment
X16361 N16361 N16362 Segment
X16362 N16362 N16363 Segment
X16363 N16363 N16364 Segment
X16364 N16364 N16365 Segment
X16365 N16365 N16366 Segment
X16366 N16366 N16367 Segment
X16367 N16367 N16368 Segment
X16368 N16368 N16369 Segment
X16369 N16369 N16370 Segment
X16370 N16370 N16371 Segment
X16371 N16371 N16372 Segment
X16372 N16372 N16373 Segment
X16373 N16373 N16374 Segment
X16374 N16374 N16375 Segment
X16375 N16375 N16376 Segment
X16376 N16376 N16377 Segment
X16377 N16377 N16378 Segment
X16378 N16378 N16379 Segment
X16379 N16379 N16380 Segment
X16380 N16380 N16381 Segment
X16381 N16381 N16382 Segment
X16382 N16382 N16383 Segment
X16383 N16383 N16384 Segment
X16384 N16384 N16385 Segment
X16385 N16385 N16386 Segment
X16386 N16386 N16387 Segment
X16387 N16387 N16388 Segment
X16388 N16388 N16389 Segment
X16389 N16389 N16390 Segment
X16390 N16390 N16391 Segment
X16391 N16391 N16392 Segment
X16392 N16392 N16393 Segment
X16393 N16393 N16394 Segment
X16394 N16394 N16395 Segment
X16395 N16395 N16396 Segment
X16396 N16396 N16397 Segment
X16397 N16397 N16398 Segment
X16398 N16398 N16399 Segment
X16399 N16399 N16400 Segment
X16400 N16400 N16401 Segment
X16401 N16401 N16402 Segment
X16402 N16402 N16403 Segment
X16403 N16403 N16404 Segment
X16404 N16404 N16405 Segment
X16405 N16405 N16406 Segment
X16406 N16406 N16407 Segment
X16407 N16407 N16408 Segment
X16408 N16408 N16409 Segment
X16409 N16409 N16410 Segment
X16410 N16410 N16411 Segment
X16411 N16411 N16412 Segment
X16412 N16412 N16413 Segment
X16413 N16413 N16414 Segment
X16414 N16414 N16415 Segment
X16415 N16415 N16416 Segment
X16416 N16416 N16417 Segment
X16417 N16417 N16418 Segment
X16418 N16418 N16419 Segment
X16419 N16419 N16420 Segment
X16420 N16420 N16421 Segment
X16421 N16421 N16422 Segment
X16422 N16422 N16423 Segment
X16423 N16423 N16424 Segment
X16424 N16424 N16425 Segment
X16425 N16425 N16426 Segment
X16426 N16426 N16427 Segment
X16427 N16427 N16428 Segment
X16428 N16428 N16429 Segment
X16429 N16429 N16430 Segment
X16430 N16430 N16431 Segment
X16431 N16431 N16432 Segment
X16432 N16432 N16433 Segment
X16433 N16433 N16434 Segment
X16434 N16434 N16435 Segment
X16435 N16435 N16436 Segment
X16436 N16436 N16437 Segment
X16437 N16437 N16438 Segment
X16438 N16438 N16439 Segment
X16439 N16439 N16440 Segment
X16440 N16440 N16441 Segment
X16441 N16441 N16442 Segment
X16442 N16442 N16443 Segment
X16443 N16443 N16444 Segment
X16444 N16444 N16445 Segment
X16445 N16445 N16446 Segment
X16446 N16446 N16447 Segment
X16447 N16447 N16448 Segment
X16448 N16448 N16449 Segment
X16449 N16449 N16450 Segment
X16450 N16450 N16451 Segment
X16451 N16451 N16452 Segment
X16452 N16452 N16453 Segment
X16453 N16453 N16454 Segment
X16454 N16454 N16455 Segment
X16455 N16455 N16456 Segment
X16456 N16456 N16457 Segment
X16457 N16457 N16458 Segment
X16458 N16458 N16459 Segment
X16459 N16459 N16460 Segment
X16460 N16460 N16461 Segment
X16461 N16461 N16462 Segment
X16462 N16462 N16463 Segment
X16463 N16463 N16464 Segment
X16464 N16464 N16465 Segment
X16465 N16465 N16466 Segment
X16466 N16466 N16467 Segment
X16467 N16467 N16468 Segment
X16468 N16468 N16469 Segment
X16469 N16469 N16470 Segment
X16470 N16470 N16471 Segment
X16471 N16471 N16472 Segment
X16472 N16472 N16473 Segment
X16473 N16473 N16474 Segment
X16474 N16474 N16475 Segment
X16475 N16475 N16476 Segment
X16476 N16476 N16477 Segment
X16477 N16477 N16478 Segment
X16478 N16478 N16479 Segment
X16479 N16479 N16480 Segment
X16480 N16480 N16481 Segment
X16481 N16481 N16482 Segment
X16482 N16482 N16483 Segment
X16483 N16483 N16484 Segment
X16484 N16484 N16485 Segment
X16485 N16485 N16486 Segment
X16486 N16486 N16487 Segment
X16487 N16487 N16488 Segment
X16488 N16488 N16489 Segment
X16489 N16489 N16490 Segment
X16490 N16490 N16491 Segment
X16491 N16491 N16492 Segment
X16492 N16492 N16493 Segment
X16493 N16493 N16494 Segment
X16494 N16494 N16495 Segment
X16495 N16495 N16496 Segment
X16496 N16496 N16497 Segment
X16497 N16497 N16498 Segment
X16498 N16498 N16499 Segment
X16499 N16499 N16500 Segment
X16500 N16500 N16501 Segment
X16501 N16501 N16502 Segment
X16502 N16502 N16503 Segment
X16503 N16503 N16504 Segment
X16504 N16504 N16505 Segment
X16505 N16505 N16506 Segment
X16506 N16506 N16507 Segment
X16507 N16507 N16508 Segment
X16508 N16508 N16509 Segment
X16509 N16509 N16510 Segment
X16510 N16510 N16511 Segment
X16511 N16511 N16512 Segment
X16512 N16512 N16513 Segment
X16513 N16513 N16514 Segment
X16514 N16514 N16515 Segment
X16515 N16515 N16516 Segment
X16516 N16516 N16517 Segment
X16517 N16517 N16518 Segment
X16518 N16518 N16519 Segment
X16519 N16519 N16520 Segment
X16520 N16520 N16521 Segment
X16521 N16521 N16522 Segment
X16522 N16522 N16523 Segment
X16523 N16523 N16524 Segment
X16524 N16524 N16525 Segment
X16525 N16525 N16526 Segment
X16526 N16526 N16527 Segment
X16527 N16527 N16528 Segment
X16528 N16528 N16529 Segment
X16529 N16529 N16530 Segment
X16530 N16530 N16531 Segment
X16531 N16531 N16532 Segment
X16532 N16532 N16533 Segment
X16533 N16533 N16534 Segment
X16534 N16534 N16535 Segment
X16535 N16535 N16536 Segment
X16536 N16536 N16537 Segment
X16537 N16537 N16538 Segment
X16538 N16538 N16539 Segment
X16539 N16539 N16540 Segment
X16540 N16540 N16541 Segment
X16541 N16541 N16542 Segment
X16542 N16542 N16543 Segment
X16543 N16543 N16544 Segment
X16544 N16544 N16545 Segment
X16545 N16545 N16546 Segment
X16546 N16546 N16547 Segment
X16547 N16547 N16548 Segment
X16548 N16548 N16549 Segment
X16549 N16549 N16550 Segment
X16550 N16550 N16551 Segment
X16551 N16551 N16552 Segment
X16552 N16552 N16553 Segment
X16553 N16553 N16554 Segment
X16554 N16554 N16555 Segment
X16555 N16555 N16556 Segment
X16556 N16556 N16557 Segment
X16557 N16557 N16558 Segment
X16558 N16558 N16559 Segment
X16559 N16559 N16560 Segment
X16560 N16560 N16561 Segment
X16561 N16561 N16562 Segment
X16562 N16562 N16563 Segment
X16563 N16563 N16564 Segment
X16564 N16564 N16565 Segment
X16565 N16565 N16566 Segment
X16566 N16566 N16567 Segment
X16567 N16567 N16568 Segment
X16568 N16568 N16569 Segment
X16569 N16569 N16570 Segment
X16570 N16570 N16571 Segment
X16571 N16571 N16572 Segment
X16572 N16572 N16573 Segment
X16573 N16573 N16574 Segment
X16574 N16574 N16575 Segment
X16575 N16575 N16576 Segment
X16576 N16576 N16577 Segment
X16577 N16577 N16578 Segment
X16578 N16578 N16579 Segment
X16579 N16579 N16580 Segment
X16580 N16580 N16581 Segment
X16581 N16581 N16582 Segment
X16582 N16582 N16583 Segment
X16583 N16583 N16584 Segment
X16584 N16584 N16585 Segment
X16585 N16585 N16586 Segment
X16586 N16586 N16587 Segment
X16587 N16587 N16588 Segment
X16588 N16588 N16589 Segment
X16589 N16589 N16590 Segment
X16590 N16590 N16591 Segment
X16591 N16591 N16592 Segment
X16592 N16592 N16593 Segment
X16593 N16593 N16594 Segment
X16594 N16594 N16595 Segment
X16595 N16595 N16596 Segment
X16596 N16596 N16597 Segment
X16597 N16597 N16598 Segment
X16598 N16598 N16599 Segment
X16599 N16599 N16600 Segment
X16600 N16600 N16601 Segment
X16601 N16601 N16602 Segment
X16602 N16602 N16603 Segment
X16603 N16603 N16604 Segment
X16604 N16604 N16605 Segment
X16605 N16605 N16606 Segment
X16606 N16606 N16607 Segment
X16607 N16607 N16608 Segment
X16608 N16608 N16609 Segment
X16609 N16609 N16610 Segment
X16610 N16610 N16611 Segment
X16611 N16611 N16612 Segment
X16612 N16612 N16613 Segment
X16613 N16613 N16614 Segment
X16614 N16614 N16615 Segment
X16615 N16615 N16616 Segment
X16616 N16616 N16617 Segment
X16617 N16617 N16618 Segment
X16618 N16618 N16619 Segment
X16619 N16619 N16620 Segment
X16620 N16620 N16621 Segment
X16621 N16621 N16622 Segment
X16622 N16622 N16623 Segment
X16623 N16623 N16624 Segment
X16624 N16624 N16625 Segment
X16625 N16625 N16626 Segment
X16626 N16626 N16627 Segment
X16627 N16627 N16628 Segment
X16628 N16628 N16629 Segment
X16629 N16629 N16630 Segment
X16630 N16630 N16631 Segment
X16631 N16631 N16632 Segment
X16632 N16632 N16633 Segment
X16633 N16633 N16634 Segment
X16634 N16634 N16635 Segment
X16635 N16635 N16636 Segment
X16636 N16636 N16637 Segment
X16637 N16637 N16638 Segment
X16638 N16638 N16639 Segment
X16639 N16639 N16640 Segment
X16640 N16640 N16641 Segment
X16641 N16641 N16642 Segment
X16642 N16642 N16643 Segment
X16643 N16643 N16644 Segment
X16644 N16644 N16645 Segment
X16645 N16645 N16646 Segment
X16646 N16646 N16647 Segment
X16647 N16647 N16648 Segment
X16648 N16648 N16649 Segment
X16649 N16649 N16650 Segment
X16650 N16650 N16651 Segment
X16651 N16651 N16652 Segment
X16652 N16652 N16653 Segment
X16653 N16653 N16654 Segment
X16654 N16654 N16655 Segment
X16655 N16655 N16656 Segment
X16656 N16656 N16657 Segment
X16657 N16657 N16658 Segment
X16658 N16658 N16659 Segment
X16659 N16659 N16660 Segment
X16660 N16660 N16661 Segment
X16661 N16661 N16662 Segment
X16662 N16662 N16663 Segment
X16663 N16663 N16664 Segment
X16664 N16664 N16665 Segment
X16665 N16665 N16666 Segment
X16666 N16666 N16667 Segment
X16667 N16667 N16668 Segment
X16668 N16668 N16669 Segment
X16669 N16669 N16670 Segment
X16670 N16670 N16671 Segment
X16671 N16671 N16672 Segment
X16672 N16672 N16673 Segment
X16673 N16673 N16674 Segment
X16674 N16674 N16675 Segment
X16675 N16675 N16676 Segment
X16676 N16676 N16677 Segment
X16677 N16677 N16678 Segment
X16678 N16678 N16679 Segment
X16679 N16679 N16680 Segment
X16680 N16680 N16681 Segment
X16681 N16681 N16682 Segment
X16682 N16682 N16683 Segment
X16683 N16683 N16684 Segment
X16684 N16684 N16685 Segment
X16685 N16685 N16686 Segment
X16686 N16686 N16687 Segment
X16687 N16687 N16688 Segment
X16688 N16688 N16689 Segment
X16689 N16689 N16690 Segment
X16690 N16690 N16691 Segment
X16691 N16691 N16692 Segment
X16692 N16692 N16693 Segment
X16693 N16693 N16694 Segment
X16694 N16694 N16695 Segment
X16695 N16695 N16696 Segment
X16696 N16696 N16697 Segment
X16697 N16697 N16698 Segment
X16698 N16698 N16699 Segment
X16699 N16699 N16700 Segment
X16700 N16700 N16701 Segment
X16701 N16701 N16702 Segment
X16702 N16702 N16703 Segment
X16703 N16703 N16704 Segment
X16704 N16704 N16705 Segment
X16705 N16705 N16706 Segment
X16706 N16706 N16707 Segment
X16707 N16707 N16708 Segment
X16708 N16708 N16709 Segment
X16709 N16709 N16710 Segment
X16710 N16710 N16711 Segment
X16711 N16711 N16712 Segment
X16712 N16712 N16713 Segment
X16713 N16713 N16714 Segment
X16714 N16714 N16715 Segment
X16715 N16715 N16716 Segment
X16716 N16716 N16717 Segment
X16717 N16717 N16718 Segment
X16718 N16718 N16719 Segment
X16719 N16719 N16720 Segment
X16720 N16720 N16721 Segment
X16721 N16721 N16722 Segment
X16722 N16722 N16723 Segment
X16723 N16723 N16724 Segment
X16724 N16724 N16725 Segment
X16725 N16725 N16726 Segment
X16726 N16726 N16727 Segment
X16727 N16727 N16728 Segment
X16728 N16728 N16729 Segment
X16729 N16729 N16730 Segment
X16730 N16730 N16731 Segment
X16731 N16731 N16732 Segment
X16732 N16732 N16733 Segment
X16733 N16733 N16734 Segment
X16734 N16734 N16735 Segment
X16735 N16735 N16736 Segment
X16736 N16736 N16737 Segment
X16737 N16737 N16738 Segment
X16738 N16738 N16739 Segment
X16739 N16739 N16740 Segment
X16740 N16740 N16741 Segment
X16741 N16741 N16742 Segment
X16742 N16742 N16743 Segment
X16743 N16743 N16744 Segment
X16744 N16744 N16745 Segment
X16745 N16745 N16746 Segment
X16746 N16746 N16747 Segment
X16747 N16747 N16748 Segment
X16748 N16748 N16749 Segment
X16749 N16749 N16750 Segment
X16750 N16750 N16751 Segment
X16751 N16751 N16752 Segment
X16752 N16752 N16753 Segment
X16753 N16753 N16754 Segment
X16754 N16754 N16755 Segment
X16755 N16755 N16756 Segment
X16756 N16756 N16757 Segment
X16757 N16757 N16758 Segment
X16758 N16758 N16759 Segment
X16759 N16759 N16760 Segment
X16760 N16760 N16761 Segment
X16761 N16761 N16762 Segment
X16762 N16762 N16763 Segment
X16763 N16763 N16764 Segment
X16764 N16764 N16765 Segment
X16765 N16765 N16766 Segment
X16766 N16766 N16767 Segment
X16767 N16767 N16768 Segment
X16768 N16768 N16769 Segment
X16769 N16769 N16770 Segment
X16770 N16770 N16771 Segment
X16771 N16771 N16772 Segment
X16772 N16772 N16773 Segment
X16773 N16773 N16774 Segment
X16774 N16774 N16775 Segment
X16775 N16775 N16776 Segment
X16776 N16776 N16777 Segment
X16777 N16777 N16778 Segment
X16778 N16778 N16779 Segment
X16779 N16779 N16780 Segment
X16780 N16780 N16781 Segment
X16781 N16781 N16782 Segment
X16782 N16782 N16783 Segment
X16783 N16783 N16784 Segment
X16784 N16784 N16785 Segment
X16785 N16785 N16786 Segment
X16786 N16786 N16787 Segment
X16787 N16787 N16788 Segment
X16788 N16788 N16789 Segment
X16789 N16789 N16790 Segment
X16790 N16790 N16791 Segment
X16791 N16791 N16792 Segment
X16792 N16792 N16793 Segment
X16793 N16793 N16794 Segment
X16794 N16794 N16795 Segment
X16795 N16795 N16796 Segment
X16796 N16796 N16797 Segment
X16797 N16797 N16798 Segment
X16798 N16798 N16799 Segment
X16799 N16799 N16800 Segment
X16800 N16800 N16801 Segment
X16801 N16801 N16802 Segment
X16802 N16802 N16803 Segment
X16803 N16803 N16804 Segment
X16804 N16804 N16805 Segment
X16805 N16805 N16806 Segment
X16806 N16806 N16807 Segment
X16807 N16807 N16808 Segment
X16808 N16808 N16809 Segment
X16809 N16809 N16810 Segment
X16810 N16810 N16811 Segment
X16811 N16811 N16812 Segment
X16812 N16812 N16813 Segment
X16813 N16813 N16814 Segment
X16814 N16814 N16815 Segment
X16815 N16815 N16816 Segment
X16816 N16816 N16817 Segment
X16817 N16817 N16818 Segment
X16818 N16818 N16819 Segment
X16819 N16819 N16820 Segment
X16820 N16820 N16821 Segment
X16821 N16821 N16822 Segment
X16822 N16822 N16823 Segment
X16823 N16823 N16824 Segment
X16824 N16824 N16825 Segment
X16825 N16825 N16826 Segment
X16826 N16826 N16827 Segment
X16827 N16827 N16828 Segment
X16828 N16828 N16829 Segment
X16829 N16829 N16830 Segment
X16830 N16830 N16831 Segment
X16831 N16831 N16832 Segment
X16832 N16832 N16833 Segment
X16833 N16833 N16834 Segment
X16834 N16834 N16835 Segment
X16835 N16835 N16836 Segment
X16836 N16836 N16837 Segment
X16837 N16837 N16838 Segment
X16838 N16838 N16839 Segment
X16839 N16839 N16840 Segment
X16840 N16840 N16841 Segment
X16841 N16841 N16842 Segment
X16842 N16842 N16843 Segment
X16843 N16843 N16844 Segment
X16844 N16844 N16845 Segment
X16845 N16845 N16846 Segment
X16846 N16846 N16847 Segment
X16847 N16847 N16848 Segment
X16848 N16848 N16849 Segment
X16849 N16849 N16850 Segment
X16850 N16850 N16851 Segment
X16851 N16851 N16852 Segment
X16852 N16852 N16853 Segment
X16853 N16853 N16854 Segment
X16854 N16854 N16855 Segment
X16855 N16855 N16856 Segment
X16856 N16856 N16857 Segment
X16857 N16857 N16858 Segment
X16858 N16858 N16859 Segment
X16859 N16859 N16860 Segment
X16860 N16860 N16861 Segment
X16861 N16861 N16862 Segment
X16862 N16862 N16863 Segment
X16863 N16863 N16864 Segment
X16864 N16864 N16865 Segment
X16865 N16865 N16866 Segment
X16866 N16866 N16867 Segment
X16867 N16867 N16868 Segment
X16868 N16868 N16869 Segment
X16869 N16869 N16870 Segment
X16870 N16870 N16871 Segment
X16871 N16871 N16872 Segment
X16872 N16872 N16873 Segment
X16873 N16873 N16874 Segment
X16874 N16874 N16875 Segment
X16875 N16875 N16876 Segment
X16876 N16876 N16877 Segment
X16877 N16877 N16878 Segment
X16878 N16878 N16879 Segment
X16879 N16879 N16880 Segment
X16880 N16880 N16881 Segment
X16881 N16881 N16882 Segment
X16882 N16882 N16883 Segment
X16883 N16883 N16884 Segment
X16884 N16884 N16885 Segment
X16885 N16885 N16886 Segment
X16886 N16886 N16887 Segment
X16887 N16887 N16888 Segment
X16888 N16888 N16889 Segment
X16889 N16889 N16890 Segment
X16890 N16890 N16891 Segment
X16891 N16891 N16892 Segment
X16892 N16892 N16893 Segment
X16893 N16893 N16894 Segment
X16894 N16894 N16895 Segment
X16895 N16895 N16896 Segment
X16896 N16896 N16897 Segment
X16897 N16897 N16898 Segment
X16898 N16898 N16899 Segment
X16899 N16899 N16900 Segment
X16900 N16900 N16901 Segment
X16901 N16901 N16902 Segment
X16902 N16902 N16903 Segment
X16903 N16903 N16904 Segment
X16904 N16904 N16905 Segment
X16905 N16905 N16906 Segment
X16906 N16906 N16907 Segment
X16907 N16907 N16908 Segment
X16908 N16908 N16909 Segment
X16909 N16909 N16910 Segment
X16910 N16910 N16911 Segment
X16911 N16911 N16912 Segment
X16912 N16912 N16913 Segment
X16913 N16913 N16914 Segment
X16914 N16914 N16915 Segment
X16915 N16915 N16916 Segment
X16916 N16916 N16917 Segment
X16917 N16917 N16918 Segment
X16918 N16918 N16919 Segment
X16919 N16919 N16920 Segment
X16920 N16920 N16921 Segment
X16921 N16921 N16922 Segment
X16922 N16922 N16923 Segment
X16923 N16923 N16924 Segment
X16924 N16924 N16925 Segment
X16925 N16925 N16926 Segment
X16926 N16926 N16927 Segment
X16927 N16927 N16928 Segment
X16928 N16928 N16929 Segment
X16929 N16929 N16930 Segment
X16930 N16930 N16931 Segment
X16931 N16931 N16932 Segment
X16932 N16932 N16933 Segment
X16933 N16933 N16934 Segment
X16934 N16934 N16935 Segment
X16935 N16935 N16936 Segment
X16936 N16936 N16937 Segment
X16937 N16937 N16938 Segment
X16938 N16938 N16939 Segment
X16939 N16939 N16940 Segment
X16940 N16940 N16941 Segment
X16941 N16941 N16942 Segment
X16942 N16942 N16943 Segment
X16943 N16943 N16944 Segment
X16944 N16944 N16945 Segment
X16945 N16945 N16946 Segment
X16946 N16946 N16947 Segment
X16947 N16947 N16948 Segment
X16948 N16948 N16949 Segment
X16949 N16949 N16950 Segment
X16950 N16950 N16951 Segment
X16951 N16951 N16952 Segment
X16952 N16952 N16953 Segment
X16953 N16953 N16954 Segment
X16954 N16954 N16955 Segment
X16955 N16955 N16956 Segment
X16956 N16956 N16957 Segment
X16957 N16957 N16958 Segment
X16958 N16958 N16959 Segment
X16959 N16959 N16960 Segment
X16960 N16960 N16961 Segment
X16961 N16961 N16962 Segment
X16962 N16962 N16963 Segment
X16963 N16963 N16964 Segment
X16964 N16964 N16965 Segment
X16965 N16965 N16966 Segment
X16966 N16966 N16967 Segment
X16967 N16967 N16968 Segment
X16968 N16968 N16969 Segment
X16969 N16969 N16970 Segment
X16970 N16970 N16971 Segment
X16971 N16971 N16972 Segment
X16972 N16972 N16973 Segment
X16973 N16973 N16974 Segment
X16974 N16974 N16975 Segment
X16975 N16975 N16976 Segment
X16976 N16976 N16977 Segment
X16977 N16977 N16978 Segment
X16978 N16978 N16979 Segment
X16979 N16979 N16980 Segment
X16980 N16980 N16981 Segment
X16981 N16981 N16982 Segment
X16982 N16982 N16983 Segment
X16983 N16983 N16984 Segment
X16984 N16984 N16985 Segment
X16985 N16985 N16986 Segment
X16986 N16986 N16987 Segment
X16987 N16987 N16988 Segment
X16988 N16988 N16989 Segment
X16989 N16989 N16990 Segment
X16990 N16990 N16991 Segment
X16991 N16991 N16992 Segment
X16992 N16992 N16993 Segment
X16993 N16993 N16994 Segment
X16994 N16994 N16995 Segment
X16995 N16995 N16996 Segment
X16996 N16996 N16997 Segment
X16997 N16997 N16998 Segment
X16998 N16998 N16999 Segment
X16999 N16999 N17000 Segment
X17000 N17000 N17001 Segment
X17001 N17001 N17002 Segment
X17002 N17002 N17003 Segment
X17003 N17003 N17004 Segment
X17004 N17004 N17005 Segment
X17005 N17005 N17006 Segment
X17006 N17006 N17007 Segment
X17007 N17007 N17008 Segment
X17008 N17008 N17009 Segment
X17009 N17009 N17010 Segment
X17010 N17010 N17011 Segment
X17011 N17011 N17012 Segment
X17012 N17012 N17013 Segment
X17013 N17013 N17014 Segment
X17014 N17014 N17015 Segment
X17015 N17015 N17016 Segment
X17016 N17016 N17017 Segment
X17017 N17017 N17018 Segment
X17018 N17018 N17019 Segment
X17019 N17019 N17020 Segment
X17020 N17020 N17021 Segment
X17021 N17021 N17022 Segment
X17022 N17022 N17023 Segment
X17023 N17023 N17024 Segment
X17024 N17024 N17025 Segment
X17025 N17025 N17026 Segment
X17026 N17026 N17027 Segment
X17027 N17027 N17028 Segment
X17028 N17028 N17029 Segment
X17029 N17029 N17030 Segment
X17030 N17030 N17031 Segment
X17031 N17031 N17032 Segment
X17032 N17032 N17033 Segment
X17033 N17033 N17034 Segment
X17034 N17034 N17035 Segment
X17035 N17035 N17036 Segment
X17036 N17036 N17037 Segment
X17037 N17037 N17038 Segment
X17038 N17038 N17039 Segment
X17039 N17039 N17040 Segment
X17040 N17040 N17041 Segment
X17041 N17041 N17042 Segment
X17042 N17042 N17043 Segment
X17043 N17043 N17044 Segment
X17044 N17044 N17045 Segment
X17045 N17045 N17046 Segment
X17046 N17046 N17047 Segment
X17047 N17047 N17048 Segment
X17048 N17048 N17049 Segment
X17049 N17049 N17050 Segment
X17050 N17050 N17051 Segment
X17051 N17051 N17052 Segment
X17052 N17052 N17053 Segment
X17053 N17053 N17054 Segment
X17054 N17054 N17055 Segment
X17055 N17055 N17056 Segment
X17056 N17056 N17057 Segment
X17057 N17057 N17058 Segment
X17058 N17058 N17059 Segment
X17059 N17059 N17060 Segment
X17060 N17060 N17061 Segment
X17061 N17061 N17062 Segment
X17062 N17062 N17063 Segment
X17063 N17063 N17064 Segment
X17064 N17064 N17065 Segment
X17065 N17065 N17066 Segment
X17066 N17066 N17067 Segment
X17067 N17067 N17068 Segment
X17068 N17068 N17069 Segment
X17069 N17069 N17070 Segment
X17070 N17070 N17071 Segment
X17071 N17071 N17072 Segment
X17072 N17072 N17073 Segment
X17073 N17073 N17074 Segment
X17074 N17074 N17075 Segment
X17075 N17075 N17076 Segment
X17076 N17076 N17077 Segment
X17077 N17077 N17078 Segment
X17078 N17078 N17079 Segment
X17079 N17079 N17080 Segment
X17080 N17080 N17081 Segment
X17081 N17081 N17082 Segment
X17082 N17082 N17083 Segment
X17083 N17083 N17084 Segment
X17084 N17084 N17085 Segment
X17085 N17085 N17086 Segment
X17086 N17086 N17087 Segment
X17087 N17087 N17088 Segment
X17088 N17088 N17089 Segment
X17089 N17089 N17090 Segment
X17090 N17090 N17091 Segment
X17091 N17091 N17092 Segment
X17092 N17092 N17093 Segment
X17093 N17093 N17094 Segment
X17094 N17094 N17095 Segment
X17095 N17095 N17096 Segment
X17096 N17096 N17097 Segment
X17097 N17097 N17098 Segment
X17098 N17098 N17099 Segment
X17099 N17099 N17100 Segment
X17100 N17100 N17101 Segment
X17101 N17101 N17102 Segment
X17102 N17102 N17103 Segment
X17103 N17103 N17104 Segment
X17104 N17104 N17105 Segment
X17105 N17105 N17106 Segment
X17106 N17106 N17107 Segment
X17107 N17107 N17108 Segment
X17108 N17108 N17109 Segment
X17109 N17109 N17110 Segment
X17110 N17110 N17111 Segment
X17111 N17111 N17112 Segment
X17112 N17112 N17113 Segment
X17113 N17113 N17114 Segment
X17114 N17114 N17115 Segment
X17115 N17115 N17116 Segment
X17116 N17116 N17117 Segment
X17117 N17117 N17118 Segment
X17118 N17118 N17119 Segment
X17119 N17119 N17120 Segment
X17120 N17120 N17121 Segment
X17121 N17121 N17122 Segment
X17122 N17122 N17123 Segment
X17123 N17123 N17124 Segment
X17124 N17124 N17125 Segment
X17125 N17125 N17126 Segment
X17126 N17126 N17127 Segment
X17127 N17127 N17128 Segment
X17128 N17128 N17129 Segment
X17129 N17129 N17130 Segment
X17130 N17130 N17131 Segment
X17131 N17131 N17132 Segment
X17132 N17132 N17133 Segment
X17133 N17133 N17134 Segment
X17134 N17134 N17135 Segment
X17135 N17135 N17136 Segment
X17136 N17136 N17137 Segment
X17137 N17137 N17138 Segment
X17138 N17138 N17139 Segment
X17139 N17139 N17140 Segment
X17140 N17140 N17141 Segment
X17141 N17141 N17142 Segment
X17142 N17142 N17143 Segment
X17143 N17143 N17144 Segment
X17144 N17144 N17145 Segment
X17145 N17145 N17146 Segment
X17146 N17146 N17147 Segment
X17147 N17147 N17148 Segment
X17148 N17148 N17149 Segment
X17149 N17149 N17150 Segment
X17150 N17150 N17151 Segment
X17151 N17151 N17152 Segment
X17152 N17152 N17153 Segment
X17153 N17153 N17154 Segment
X17154 N17154 N17155 Segment
X17155 N17155 N17156 Segment
X17156 N17156 N17157 Segment
X17157 N17157 N17158 Segment
X17158 N17158 N17159 Segment
X17159 N17159 N17160 Segment
X17160 N17160 N17161 Segment
X17161 N17161 N17162 Segment
X17162 N17162 N17163 Segment
X17163 N17163 N17164 Segment
X17164 N17164 N17165 Segment
X17165 N17165 N17166 Segment
X17166 N17166 N17167 Segment
X17167 N17167 N17168 Segment
X17168 N17168 N17169 Segment
X17169 N17169 N17170 Segment
X17170 N17170 N17171 Segment
X17171 N17171 N17172 Segment
X17172 N17172 N17173 Segment
X17173 N17173 N17174 Segment
X17174 N17174 N17175 Segment
X17175 N17175 N17176 Segment
X17176 N17176 N17177 Segment
X17177 N17177 N17178 Segment
X17178 N17178 N17179 Segment
X17179 N17179 N17180 Segment
X17180 N17180 N17181 Segment
X17181 N17181 N17182 Segment
X17182 N17182 N17183 Segment
X17183 N17183 N17184 Segment
X17184 N17184 N17185 Segment
X17185 N17185 N17186 Segment
X17186 N17186 N17187 Segment
X17187 N17187 N17188 Segment
X17188 N17188 N17189 Segment
X17189 N17189 N17190 Segment
X17190 N17190 N17191 Segment
X17191 N17191 N17192 Segment
X17192 N17192 N17193 Segment
X17193 N17193 N17194 Segment
X17194 N17194 N17195 Segment
X17195 N17195 N17196 Segment
X17196 N17196 N17197 Segment
X17197 N17197 N17198 Segment
X17198 N17198 N17199 Segment
X17199 N17199 N17200 Segment
X17200 N17200 N17201 Segment
X17201 N17201 N17202 Segment
X17202 N17202 N17203 Segment
X17203 N17203 N17204 Segment
X17204 N17204 N17205 Segment
X17205 N17205 N17206 Segment
X17206 N17206 N17207 Segment
X17207 N17207 N17208 Segment
X17208 N17208 N17209 Segment
X17209 N17209 N17210 Segment
X17210 N17210 N17211 Segment
X17211 N17211 N17212 Segment
X17212 N17212 N17213 Segment
X17213 N17213 N17214 Segment
X17214 N17214 N17215 Segment
X17215 N17215 N17216 Segment
X17216 N17216 N17217 Segment
X17217 N17217 N17218 Segment
X17218 N17218 N17219 Segment
X17219 N17219 N17220 Segment
X17220 N17220 N17221 Segment
X17221 N17221 N17222 Segment
X17222 N17222 N17223 Segment
X17223 N17223 N17224 Segment
X17224 N17224 N17225 Segment
X17225 N17225 N17226 Segment
X17226 N17226 N17227 Segment
X17227 N17227 N17228 Segment
X17228 N17228 N17229 Segment
X17229 N17229 N17230 Segment
X17230 N17230 N17231 Segment
X17231 N17231 N17232 Segment
X17232 N17232 N17233 Segment
X17233 N17233 N17234 Segment
X17234 N17234 N17235 Segment
X17235 N17235 N17236 Segment
X17236 N17236 N17237 Segment
X17237 N17237 N17238 Segment
X17238 N17238 N17239 Segment
X17239 N17239 N17240 Segment
X17240 N17240 N17241 Segment
X17241 N17241 N17242 Segment
X17242 N17242 N17243 Segment
X17243 N17243 N17244 Segment
X17244 N17244 N17245 Segment
X17245 N17245 N17246 Segment
X17246 N17246 N17247 Segment
X17247 N17247 N17248 Segment
X17248 N17248 N17249 Segment
X17249 N17249 N17250 Segment
X17250 N17250 N17251 Segment
X17251 N17251 N17252 Segment
X17252 N17252 N17253 Segment
X17253 N17253 N17254 Segment
X17254 N17254 N17255 Segment
X17255 N17255 N17256 Segment
X17256 N17256 N17257 Segment
X17257 N17257 N17258 Segment
X17258 N17258 N17259 Segment
X17259 N17259 N17260 Segment
X17260 N17260 N17261 Segment
X17261 N17261 N17262 Segment
X17262 N17262 N17263 Segment
X17263 N17263 N17264 Segment
X17264 N17264 N17265 Segment
X17265 N17265 N17266 Segment
X17266 N17266 N17267 Segment
X17267 N17267 N17268 Segment
X17268 N17268 N17269 Segment
X17269 N17269 N17270 Segment
X17270 N17270 N17271 Segment
X17271 N17271 N17272 Segment
X17272 N17272 N17273 Segment
X17273 N17273 N17274 Segment
X17274 N17274 N17275 Segment
X17275 N17275 N17276 Segment
X17276 N17276 N17277 Segment
X17277 N17277 N17278 Segment
X17278 N17278 N17279 Segment
X17279 N17279 N17280 Segment
X17280 N17280 N17281 Segment
X17281 N17281 N17282 Segment
X17282 N17282 N17283 Segment
X17283 N17283 N17284 Segment
X17284 N17284 N17285 Segment
X17285 N17285 N17286 Segment
X17286 N17286 N17287 Segment
X17287 N17287 N17288 Segment
X17288 N17288 N17289 Segment
X17289 N17289 N17290 Segment
X17290 N17290 N17291 Segment
X17291 N17291 N17292 Segment
X17292 N17292 N17293 Segment
X17293 N17293 N17294 Segment
X17294 N17294 N17295 Segment
X17295 N17295 N17296 Segment
X17296 N17296 N17297 Segment
X17297 N17297 N17298 Segment
X17298 N17298 N17299 Segment
X17299 N17299 N17300 Segment
X17300 N17300 N17301 Segment
X17301 N17301 N17302 Segment
X17302 N17302 N17303 Segment
X17303 N17303 N17304 Segment
X17304 N17304 N17305 Segment
X17305 N17305 N17306 Segment
X17306 N17306 N17307 Segment
X17307 N17307 N17308 Segment
X17308 N17308 N17309 Segment
X17309 N17309 N17310 Segment
X17310 N17310 N17311 Segment
X17311 N17311 N17312 Segment
X17312 N17312 N17313 Segment
X17313 N17313 N17314 Segment
X17314 N17314 N17315 Segment
X17315 N17315 N17316 Segment
X17316 N17316 N17317 Segment
X17317 N17317 N17318 Segment
X17318 N17318 N17319 Segment
X17319 N17319 N17320 Segment
X17320 N17320 N17321 Segment
X17321 N17321 N17322 Segment
X17322 N17322 N17323 Segment
X17323 N17323 N17324 Segment
X17324 N17324 N17325 Segment
X17325 N17325 N17326 Segment
X17326 N17326 N17327 Segment
X17327 N17327 N17328 Segment
X17328 N17328 N17329 Segment
X17329 N17329 N17330 Segment
X17330 N17330 N17331 Segment
X17331 N17331 N17332 Segment
X17332 N17332 N17333 Segment
X17333 N17333 N17334 Segment
X17334 N17334 N17335 Segment
X17335 N17335 N17336 Segment
X17336 N17336 N17337 Segment
X17337 N17337 N17338 Segment
X17338 N17338 N17339 Segment
X17339 N17339 N17340 Segment
X17340 N17340 N17341 Segment
X17341 N17341 N17342 Segment
X17342 N17342 N17343 Segment
X17343 N17343 N17344 Segment
X17344 N17344 N17345 Segment
X17345 N17345 N17346 Segment
X17346 N17346 N17347 Segment
X17347 N17347 N17348 Segment
X17348 N17348 N17349 Segment
X17349 N17349 N17350 Segment
X17350 N17350 N17351 Segment
X17351 N17351 N17352 Segment
X17352 N17352 N17353 Segment
X17353 N17353 N17354 Segment
X17354 N17354 N17355 Segment
X17355 N17355 N17356 Segment
X17356 N17356 N17357 Segment
X17357 N17357 N17358 Segment
X17358 N17358 N17359 Segment
X17359 N17359 N17360 Segment
X17360 N17360 N17361 Segment
X17361 N17361 N17362 Segment
X17362 N17362 N17363 Segment
X17363 N17363 N17364 Segment
X17364 N17364 N17365 Segment
X17365 N17365 N17366 Segment
X17366 N17366 N17367 Segment
X17367 N17367 N17368 Segment
X17368 N17368 N17369 Segment
X17369 N17369 N17370 Segment
X17370 N17370 N17371 Segment
X17371 N17371 N17372 Segment
X17372 N17372 N17373 Segment
X17373 N17373 N17374 Segment
X17374 N17374 N17375 Segment
X17375 N17375 N17376 Segment
X17376 N17376 N17377 Segment
X17377 N17377 N17378 Segment
X17378 N17378 N17379 Segment
X17379 N17379 N17380 Segment
X17380 N17380 N17381 Segment
X17381 N17381 N17382 Segment
X17382 N17382 N17383 Segment
X17383 N17383 N17384 Segment
X17384 N17384 N17385 Segment
X17385 N17385 N17386 Segment
X17386 N17386 N17387 Segment
X17387 N17387 N17388 Segment
X17388 N17388 N17389 Segment
X17389 N17389 N17390 Segment
X17390 N17390 N17391 Segment
X17391 N17391 N17392 Segment
X17392 N17392 N17393 Segment
X17393 N17393 N17394 Segment
X17394 N17394 N17395 Segment
X17395 N17395 N17396 Segment
X17396 N17396 N17397 Segment
X17397 N17397 N17398 Segment
X17398 N17398 N17399 Segment
X17399 N17399 N17400 Segment
X17400 N17400 N17401 Segment
X17401 N17401 N17402 Segment
X17402 N17402 N17403 Segment
X17403 N17403 N17404 Segment
X17404 N17404 N17405 Segment
X17405 N17405 N17406 Segment
X17406 N17406 N17407 Segment
X17407 N17407 N17408 Segment
X17408 N17408 N17409 Segment
X17409 N17409 N17410 Segment
X17410 N17410 N17411 Segment
X17411 N17411 N17412 Segment
X17412 N17412 N17413 Segment
X17413 N17413 N17414 Segment
X17414 N17414 N17415 Segment
X17415 N17415 N17416 Segment
X17416 N17416 N17417 Segment
X17417 N17417 N17418 Segment
X17418 N17418 N17419 Segment
X17419 N17419 N17420 Segment
X17420 N17420 N17421 Segment
X17421 N17421 N17422 Segment
X17422 N17422 N17423 Segment
X17423 N17423 N17424 Segment
X17424 N17424 N17425 Segment
X17425 N17425 N17426 Segment
X17426 N17426 N17427 Segment
X17427 N17427 N17428 Segment
X17428 N17428 N17429 Segment
X17429 N17429 N17430 Segment
X17430 N17430 N17431 Segment
X17431 N17431 N17432 Segment
X17432 N17432 N17433 Segment
X17433 N17433 N17434 Segment
X17434 N17434 N17435 Segment
X17435 N17435 N17436 Segment
X17436 N17436 N17437 Segment
X17437 N17437 N17438 Segment
X17438 N17438 N17439 Segment
X17439 N17439 N17440 Segment
X17440 N17440 N17441 Segment
X17441 N17441 N17442 Segment
X17442 N17442 N17443 Segment
X17443 N17443 N17444 Segment
X17444 N17444 N17445 Segment
X17445 N17445 N17446 Segment
X17446 N17446 N17447 Segment
X17447 N17447 N17448 Segment
X17448 N17448 N17449 Segment
X17449 N17449 N17450 Segment
X17450 N17450 N17451 Segment
X17451 N17451 N17452 Segment
X17452 N17452 N17453 Segment
X17453 N17453 N17454 Segment
X17454 N17454 N17455 Segment
X17455 N17455 N17456 Segment
X17456 N17456 N17457 Segment
X17457 N17457 N17458 Segment
X17458 N17458 N17459 Segment
X17459 N17459 N17460 Segment
X17460 N17460 N17461 Segment
X17461 N17461 N17462 Segment
X17462 N17462 N17463 Segment
X17463 N17463 N17464 Segment
X17464 N17464 N17465 Segment
X17465 N17465 N17466 Segment
X17466 N17466 N17467 Segment
X17467 N17467 N17468 Segment
X17468 N17468 N17469 Segment
X17469 N17469 N17470 Segment
X17470 N17470 N17471 Segment
X17471 N17471 N17472 Segment
X17472 N17472 N17473 Segment
X17473 N17473 N17474 Segment
X17474 N17474 N17475 Segment
X17475 N17475 N17476 Segment
X17476 N17476 N17477 Segment
X17477 N17477 N17478 Segment
X17478 N17478 N17479 Segment
X17479 N17479 N17480 Segment
X17480 N17480 N17481 Segment
X17481 N17481 N17482 Segment
X17482 N17482 N17483 Segment
X17483 N17483 N17484 Segment
X17484 N17484 N17485 Segment
X17485 N17485 N17486 Segment
X17486 N17486 N17487 Segment
X17487 N17487 N17488 Segment
X17488 N17488 N17489 Segment
X17489 N17489 N17490 Segment
X17490 N17490 N17491 Segment
X17491 N17491 N17492 Segment
X17492 N17492 N17493 Segment
X17493 N17493 N17494 Segment
X17494 N17494 N17495 Segment
X17495 N17495 N17496 Segment
X17496 N17496 N17497 Segment
X17497 N17497 N17498 Segment
X17498 N17498 N17499 Segment
X17499 N17499 N17500 Segment
X17500 N17500 N17501 Segment
X17501 N17501 N17502 Segment
X17502 N17502 N17503 Segment
X17503 N17503 N17504 Segment
X17504 N17504 N17505 Segment
X17505 N17505 N17506 Segment
X17506 N17506 N17507 Segment
X17507 N17507 N17508 Segment
X17508 N17508 N17509 Segment
X17509 N17509 N17510 Segment
X17510 N17510 N17511 Segment
X17511 N17511 N17512 Segment
X17512 N17512 N17513 Segment
X17513 N17513 N17514 Segment
X17514 N17514 N17515 Segment
X17515 N17515 N17516 Segment
X17516 N17516 N17517 Segment
X17517 N17517 N17518 Segment
X17518 N17518 N17519 Segment
X17519 N17519 N17520 Segment
X17520 N17520 N17521 Segment
X17521 N17521 N17522 Segment
X17522 N17522 N17523 Segment
X17523 N17523 N17524 Segment
X17524 N17524 N17525 Segment
X17525 N17525 N17526 Segment
X17526 N17526 N17527 Segment
X17527 N17527 N17528 Segment
X17528 N17528 N17529 Segment
X17529 N17529 N17530 Segment
X17530 N17530 N17531 Segment
X17531 N17531 N17532 Segment
X17532 N17532 N17533 Segment
X17533 N17533 N17534 Segment
X17534 N17534 N17535 Segment
X17535 N17535 N17536 Segment
X17536 N17536 N17537 Segment
X17537 N17537 N17538 Segment
X17538 N17538 N17539 Segment
X17539 N17539 N17540 Segment
X17540 N17540 N17541 Segment
X17541 N17541 N17542 Segment
X17542 N17542 N17543 Segment
X17543 N17543 N17544 Segment
X17544 N17544 N17545 Segment
X17545 N17545 N17546 Segment
X17546 N17546 N17547 Segment
X17547 N17547 N17548 Segment
X17548 N17548 N17549 Segment
X17549 N17549 N17550 Segment
X17550 N17550 N17551 Segment
X17551 N17551 N17552 Segment
X17552 N17552 N17553 Segment
X17553 N17553 N17554 Segment
X17554 N17554 N17555 Segment
X17555 N17555 N17556 Segment
X17556 N17556 N17557 Segment
X17557 N17557 N17558 Segment
X17558 N17558 N17559 Segment
X17559 N17559 N17560 Segment
X17560 N17560 N17561 Segment
X17561 N17561 N17562 Segment
X17562 N17562 N17563 Segment
X17563 N17563 N17564 Segment
X17564 N17564 N17565 Segment
X17565 N17565 N17566 Segment
X17566 N17566 N17567 Segment
X17567 N17567 N17568 Segment
X17568 N17568 N17569 Segment
X17569 N17569 N17570 Segment
X17570 N17570 N17571 Segment
X17571 N17571 N17572 Segment
X17572 N17572 N17573 Segment
X17573 N17573 N17574 Segment
X17574 N17574 N17575 Segment
X17575 N17575 N17576 Segment
X17576 N17576 N17577 Segment
X17577 N17577 N17578 Segment
X17578 N17578 N17579 Segment
X17579 N17579 N17580 Segment
X17580 N17580 N17581 Segment
X17581 N17581 N17582 Segment
X17582 N17582 N17583 Segment
X17583 N17583 N17584 Segment
X17584 N17584 N17585 Segment
X17585 N17585 N17586 Segment
X17586 N17586 N17587 Segment
X17587 N17587 N17588 Segment
X17588 N17588 N17589 Segment
X17589 N17589 N17590 Segment
X17590 N17590 N17591 Segment
X17591 N17591 N17592 Segment
X17592 N17592 N17593 Segment
X17593 N17593 N17594 Segment
X17594 N17594 N17595 Segment
X17595 N17595 N17596 Segment
X17596 N17596 N17597 Segment
X17597 N17597 N17598 Segment
X17598 N17598 N17599 Segment
X17599 N17599 N17600 Segment
X17600 N17600 N17601 Segment
X17601 N17601 N17602 Segment
X17602 N17602 N17603 Segment
X17603 N17603 N17604 Segment
X17604 N17604 N17605 Segment
X17605 N17605 N17606 Segment
X17606 N17606 N17607 Segment
X17607 N17607 N17608 Segment
X17608 N17608 N17609 Segment
X17609 N17609 N17610 Segment
X17610 N17610 N17611 Segment
X17611 N17611 N17612 Segment
X17612 N17612 N17613 Segment
X17613 N17613 N17614 Segment
X17614 N17614 N17615 Segment
X17615 N17615 N17616 Segment
X17616 N17616 N17617 Segment
X17617 N17617 N17618 Segment
X17618 N17618 N17619 Segment
X17619 N17619 N17620 Segment
X17620 N17620 N17621 Segment
X17621 N17621 N17622 Segment
X17622 N17622 N17623 Segment
X17623 N17623 N17624 Segment
X17624 N17624 N17625 Segment
X17625 N17625 N17626 Segment
X17626 N17626 N17627 Segment
X17627 N17627 N17628 Segment
X17628 N17628 N17629 Segment
X17629 N17629 N17630 Segment
X17630 N17630 N17631 Segment
X17631 N17631 N17632 Segment
X17632 N17632 N17633 Segment
X17633 N17633 N17634 Segment
X17634 N17634 N17635 Segment
X17635 N17635 N17636 Segment
X17636 N17636 N17637 Segment
X17637 N17637 N17638 Segment
X17638 N17638 N17639 Segment
X17639 N17639 N17640 Segment
X17640 N17640 N17641 Segment
X17641 N17641 N17642 Segment
X17642 N17642 N17643 Segment
X17643 N17643 N17644 Segment
X17644 N17644 N17645 Segment
X17645 N17645 N17646 Segment
X17646 N17646 N17647 Segment
X17647 N17647 N17648 Segment
X17648 N17648 N17649 Segment
X17649 N17649 N17650 Segment
X17650 N17650 N17651 Segment
X17651 N17651 N17652 Segment
X17652 N17652 N17653 Segment
X17653 N17653 N17654 Segment
X17654 N17654 N17655 Segment
X17655 N17655 N17656 Segment
X17656 N17656 N17657 Segment
X17657 N17657 N17658 Segment
X17658 N17658 N17659 Segment
X17659 N17659 N17660 Segment
X17660 N17660 N17661 Segment
X17661 N17661 N17662 Segment
X17662 N17662 N17663 Segment
X17663 N17663 N17664 Segment
X17664 N17664 N17665 Segment
X17665 N17665 N17666 Segment
X17666 N17666 N17667 Segment
X17667 N17667 N17668 Segment
X17668 N17668 N17669 Segment
X17669 N17669 N17670 Segment
X17670 N17670 N17671 Segment
X17671 N17671 N17672 Segment
X17672 N17672 N17673 Segment
X17673 N17673 N17674 Segment
X17674 N17674 N17675 Segment
X17675 N17675 N17676 Segment
X17676 N17676 N17677 Segment
X17677 N17677 N17678 Segment
X17678 N17678 N17679 Segment
X17679 N17679 N17680 Segment
X17680 N17680 N17681 Segment
X17681 N17681 N17682 Segment
X17682 N17682 N17683 Segment
X17683 N17683 N17684 Segment
X17684 N17684 N17685 Segment
X17685 N17685 N17686 Segment
X17686 N17686 N17687 Segment
X17687 N17687 N17688 Segment
X17688 N17688 N17689 Segment
X17689 N17689 N17690 Segment
X17690 N17690 N17691 Segment
X17691 N17691 N17692 Segment
X17692 N17692 N17693 Segment
X17693 N17693 N17694 Segment
X17694 N17694 N17695 Segment
X17695 N17695 N17696 Segment
X17696 N17696 N17697 Segment
X17697 N17697 N17698 Segment
X17698 N17698 N17699 Segment
X17699 N17699 N17700 Segment
X17700 N17700 N17701 Segment
X17701 N17701 N17702 Segment
X17702 N17702 N17703 Segment
X17703 N17703 N17704 Segment
X17704 N17704 N17705 Segment
X17705 N17705 N17706 Segment
X17706 N17706 N17707 Segment
X17707 N17707 N17708 Segment
X17708 N17708 N17709 Segment
X17709 N17709 N17710 Segment
X17710 N17710 N17711 Segment
X17711 N17711 N17712 Segment
X17712 N17712 N17713 Segment
X17713 N17713 N17714 Segment
X17714 N17714 N17715 Segment
X17715 N17715 N17716 Segment
X17716 N17716 N17717 Segment
X17717 N17717 N17718 Segment
X17718 N17718 N17719 Segment
X17719 N17719 N17720 Segment
X17720 N17720 N17721 Segment
X17721 N17721 N17722 Segment
X17722 N17722 N17723 Segment
X17723 N17723 N17724 Segment
X17724 N17724 N17725 Segment
X17725 N17725 N17726 Segment
X17726 N17726 N17727 Segment
X17727 N17727 N17728 Segment
X17728 N17728 N17729 Segment
X17729 N17729 N17730 Segment
X17730 N17730 N17731 Segment
X17731 N17731 N17732 Segment
X17732 N17732 N17733 Segment
X17733 N17733 N17734 Segment
X17734 N17734 N17735 Segment
X17735 N17735 N17736 Segment
X17736 N17736 N17737 Segment
X17737 N17737 N17738 Segment
X17738 N17738 N17739 Segment
X17739 N17739 N17740 Segment
X17740 N17740 N17741 Segment
X17741 N17741 N17742 Segment
X17742 N17742 N17743 Segment
X17743 N17743 N17744 Segment
X17744 N17744 N17745 Segment
X17745 N17745 N17746 Segment
X17746 N17746 N17747 Segment
X17747 N17747 N17748 Segment
X17748 N17748 N17749 Segment
X17749 N17749 N17750 Segment
X17750 N17750 N17751 Segment
X17751 N17751 N17752 Segment
X17752 N17752 N17753 Segment
X17753 N17753 N17754 Segment
X17754 N17754 N17755 Segment
X17755 N17755 N17756 Segment
X17756 N17756 N17757 Segment
X17757 N17757 N17758 Segment
X17758 N17758 N17759 Segment
X17759 N17759 N17760 Segment
X17760 N17760 N17761 Segment
X17761 N17761 N17762 Segment
X17762 N17762 N17763 Segment
X17763 N17763 N17764 Segment
X17764 N17764 N17765 Segment
X17765 N17765 N17766 Segment
X17766 N17766 N17767 Segment
X17767 N17767 N17768 Segment
X17768 N17768 N17769 Segment
X17769 N17769 N17770 Segment
X17770 N17770 N17771 Segment
X17771 N17771 N17772 Segment
X17772 N17772 N17773 Segment
X17773 N17773 N17774 Segment
X17774 N17774 N17775 Segment
X17775 N17775 N17776 Segment
X17776 N17776 N17777 Segment
X17777 N17777 N17778 Segment
X17778 N17778 N17779 Segment
X17779 N17779 N17780 Segment
X17780 N17780 N17781 Segment
X17781 N17781 N17782 Segment
X17782 N17782 N17783 Segment
X17783 N17783 N17784 Segment
X17784 N17784 N17785 Segment
X17785 N17785 N17786 Segment
X17786 N17786 N17787 Segment
X17787 N17787 N17788 Segment
X17788 N17788 N17789 Segment
X17789 N17789 N17790 Segment
X17790 N17790 N17791 Segment
X17791 N17791 N17792 Segment
X17792 N17792 N17793 Segment
X17793 N17793 N17794 Segment
X17794 N17794 N17795 Segment
X17795 N17795 N17796 Segment
X17796 N17796 N17797 Segment
X17797 N17797 N17798 Segment
X17798 N17798 N17799 Segment
X17799 N17799 N17800 Segment
X17800 N17800 N17801 Segment
X17801 N17801 N17802 Segment
X17802 N17802 N17803 Segment
X17803 N17803 N17804 Segment
X17804 N17804 N17805 Segment
X17805 N17805 N17806 Segment
X17806 N17806 N17807 Segment
X17807 N17807 N17808 Segment
X17808 N17808 N17809 Segment
X17809 N17809 N17810 Segment
X17810 N17810 N17811 Segment
X17811 N17811 N17812 Segment
X17812 N17812 N17813 Segment
X17813 N17813 N17814 Segment
X17814 N17814 N17815 Segment
X17815 N17815 N17816 Segment
X17816 N17816 N17817 Segment
X17817 N17817 N17818 Segment
X17818 N17818 N17819 Segment
X17819 N17819 N17820 Segment
X17820 N17820 N17821 Segment
X17821 N17821 N17822 Segment
X17822 N17822 N17823 Segment
X17823 N17823 N17824 Segment
X17824 N17824 N17825 Segment
X17825 N17825 N17826 Segment
X17826 N17826 N17827 Segment
X17827 N17827 N17828 Segment
X17828 N17828 N17829 Segment
X17829 N17829 N17830 Segment
X17830 N17830 N17831 Segment
X17831 N17831 N17832 Segment
X17832 N17832 N17833 Segment
X17833 N17833 N17834 Segment
X17834 N17834 N17835 Segment
X17835 N17835 N17836 Segment
X17836 N17836 N17837 Segment
X17837 N17837 N17838 Segment
X17838 N17838 N17839 Segment
X17839 N17839 N17840 Segment
X17840 N17840 N17841 Segment
X17841 N17841 N17842 Segment
X17842 N17842 N17843 Segment
X17843 N17843 N17844 Segment
X17844 N17844 N17845 Segment
X17845 N17845 N17846 Segment
X17846 N17846 N17847 Segment
X17847 N17847 N17848 Segment
X17848 N17848 N17849 Segment
X17849 N17849 N17850 Segment
X17850 N17850 N17851 Segment
X17851 N17851 N17852 Segment
X17852 N17852 N17853 Segment
X17853 N17853 N17854 Segment
X17854 N17854 N17855 Segment
X17855 N17855 N17856 Segment
X17856 N17856 N17857 Segment
X17857 N17857 N17858 Segment
X17858 N17858 N17859 Segment
X17859 N17859 N17860 Segment
X17860 N17860 N17861 Segment
X17861 N17861 N17862 Segment
X17862 N17862 N17863 Segment
X17863 N17863 N17864 Segment
X17864 N17864 N17865 Segment
X17865 N17865 N17866 Segment
X17866 N17866 N17867 Segment
X17867 N17867 N17868 Segment
X17868 N17868 N17869 Segment
X17869 N17869 N17870 Segment
X17870 N17870 N17871 Segment
X17871 N17871 N17872 Segment
X17872 N17872 N17873 Segment
X17873 N17873 N17874 Segment
X17874 N17874 N17875 Segment
X17875 N17875 N17876 Segment
X17876 N17876 N17877 Segment
X17877 N17877 N17878 Segment
X17878 N17878 N17879 Segment
X17879 N17879 N17880 Segment
X17880 N17880 N17881 Segment
X17881 N17881 N17882 Segment
X17882 N17882 N17883 Segment
X17883 N17883 N17884 Segment
X17884 N17884 N17885 Segment
X17885 N17885 N17886 Segment
X17886 N17886 N17887 Segment
X17887 N17887 N17888 Segment
X17888 N17888 N17889 Segment
X17889 N17889 N17890 Segment
X17890 N17890 N17891 Segment
X17891 N17891 N17892 Segment
X17892 N17892 N17893 Segment
X17893 N17893 N17894 Segment
X17894 N17894 N17895 Segment
X17895 N17895 N17896 Segment
X17896 N17896 N17897 Segment
X17897 N17897 N17898 Segment
X17898 N17898 N17899 Segment
X17899 N17899 N17900 Segment
X17900 N17900 N17901 Segment
X17901 N17901 N17902 Segment
X17902 N17902 N17903 Segment
X17903 N17903 N17904 Segment
X17904 N17904 N17905 Segment
X17905 N17905 N17906 Segment
X17906 N17906 N17907 Segment
X17907 N17907 N17908 Segment
X17908 N17908 N17909 Segment
X17909 N17909 N17910 Segment
X17910 N17910 N17911 Segment
X17911 N17911 N17912 Segment
X17912 N17912 N17913 Segment
X17913 N17913 N17914 Segment
X17914 N17914 N17915 Segment
X17915 N17915 N17916 Segment
X17916 N17916 N17917 Segment
X17917 N17917 N17918 Segment
X17918 N17918 N17919 Segment
X17919 N17919 N17920 Segment
X17920 N17920 N17921 Segment
X17921 N17921 N17922 Segment
X17922 N17922 N17923 Segment
X17923 N17923 N17924 Segment
X17924 N17924 N17925 Segment
X17925 N17925 N17926 Segment
X17926 N17926 N17927 Segment
X17927 N17927 N17928 Segment
X17928 N17928 N17929 Segment
X17929 N17929 N17930 Segment
X17930 N17930 N17931 Segment
X17931 N17931 N17932 Segment
X17932 N17932 N17933 Segment
X17933 N17933 N17934 Segment
X17934 N17934 N17935 Segment
X17935 N17935 N17936 Segment
X17936 N17936 N17937 Segment
X17937 N17937 N17938 Segment
X17938 N17938 N17939 Segment
X17939 N17939 N17940 Segment
X17940 N17940 N17941 Segment
X17941 N17941 N17942 Segment
X17942 N17942 N17943 Segment
X17943 N17943 N17944 Segment
X17944 N17944 N17945 Segment
X17945 N17945 N17946 Segment
X17946 N17946 N17947 Segment
X17947 N17947 N17948 Segment
X17948 N17948 N17949 Segment
X17949 N17949 N17950 Segment
X17950 N17950 N17951 Segment
X17951 N17951 N17952 Segment
X17952 N17952 N17953 Segment
X17953 N17953 N17954 Segment
X17954 N17954 N17955 Segment
X17955 N17955 N17956 Segment
X17956 N17956 N17957 Segment
X17957 N17957 N17958 Segment
X17958 N17958 N17959 Segment
X17959 N17959 N17960 Segment
X17960 N17960 N17961 Segment
X17961 N17961 N17962 Segment
X17962 N17962 N17963 Segment
X17963 N17963 N17964 Segment
X17964 N17964 N17965 Segment
X17965 N17965 N17966 Segment
X17966 N17966 N17967 Segment
X17967 N17967 N17968 Segment
X17968 N17968 N17969 Segment
X17969 N17969 N17970 Segment
X17970 N17970 N17971 Segment
X17971 N17971 N17972 Segment
X17972 N17972 N17973 Segment
X17973 N17973 N17974 Segment
X17974 N17974 N17975 Segment
X17975 N17975 N17976 Segment
X17976 N17976 N17977 Segment
X17977 N17977 N17978 Segment
X17978 N17978 N17979 Segment
X17979 N17979 N17980 Segment
X17980 N17980 N17981 Segment
X17981 N17981 N17982 Segment
X17982 N17982 N17983 Segment
X17983 N17983 N17984 Segment
X17984 N17984 N17985 Segment
X17985 N17985 N17986 Segment
X17986 N17986 N17987 Segment
X17987 N17987 N17988 Segment
X17988 N17988 N17989 Segment
X17989 N17989 N17990 Segment
X17990 N17990 N17991 Segment
X17991 N17991 N17992 Segment
X17992 N17992 N17993 Segment
X17993 N17993 N17994 Segment
X17994 N17994 N17995 Segment
X17995 N17995 N17996 Segment
X17996 N17996 N17997 Segment
X17997 N17997 N17998 Segment
X17998 N17998 N17999 Segment
X17999 N17999 N18000 Segment
X18000 N18000 N18001 Segment
X18001 N18001 N18002 Segment
X18002 N18002 N18003 Segment
X18003 N18003 N18004 Segment
X18004 N18004 N18005 Segment
X18005 N18005 N18006 Segment
X18006 N18006 N18007 Segment
X18007 N18007 N18008 Segment
X18008 N18008 N18009 Segment
X18009 N18009 N18010 Segment
X18010 N18010 N18011 Segment
X18011 N18011 N18012 Segment
X18012 N18012 N18013 Segment
X18013 N18013 N18014 Segment
X18014 N18014 N18015 Segment
X18015 N18015 N18016 Segment
X18016 N18016 N18017 Segment
X18017 N18017 N18018 Segment
X18018 N18018 N18019 Segment
X18019 N18019 N18020 Segment
X18020 N18020 N18021 Segment
X18021 N18021 N18022 Segment
X18022 N18022 N18023 Segment
X18023 N18023 N18024 Segment
X18024 N18024 N18025 Segment
X18025 N18025 N18026 Segment
X18026 N18026 N18027 Segment
X18027 N18027 N18028 Segment
X18028 N18028 N18029 Segment
X18029 N18029 N18030 Segment
X18030 N18030 N18031 Segment
X18031 N18031 N18032 Segment
X18032 N18032 N18033 Segment
X18033 N18033 N18034 Segment
X18034 N18034 N18035 Segment
X18035 N18035 N18036 Segment
X18036 N18036 N18037 Segment
X18037 N18037 N18038 Segment
X18038 N18038 N18039 Segment
X18039 N18039 N18040 Segment
X18040 N18040 N18041 Segment
X18041 N18041 N18042 Segment
X18042 N18042 N18043 Segment
X18043 N18043 N18044 Segment
X18044 N18044 N18045 Segment
X18045 N18045 N18046 Segment
X18046 N18046 N18047 Segment
X18047 N18047 N18048 Segment
X18048 N18048 N18049 Segment
X18049 N18049 N18050 Segment
X18050 N18050 N18051 Segment
X18051 N18051 N18052 Segment
X18052 N18052 N18053 Segment
X18053 N18053 N18054 Segment
X18054 N18054 N18055 Segment
X18055 N18055 N18056 Segment
X18056 N18056 N18057 Segment
X18057 N18057 N18058 Segment
X18058 N18058 N18059 Segment
X18059 N18059 N18060 Segment
X18060 N18060 N18061 Segment
X18061 N18061 N18062 Segment
X18062 N18062 N18063 Segment
X18063 N18063 N18064 Segment
X18064 N18064 N18065 Segment
X18065 N18065 N18066 Segment
X18066 N18066 N18067 Segment
X18067 N18067 N18068 Segment
X18068 N18068 N18069 Segment
X18069 N18069 N18070 Segment
X18070 N18070 N18071 Segment
X18071 N18071 N18072 Segment
X18072 N18072 N18073 Segment
X18073 N18073 N18074 Segment
X18074 N18074 N18075 Segment
X18075 N18075 N18076 Segment
X18076 N18076 N18077 Segment
X18077 N18077 N18078 Segment
X18078 N18078 N18079 Segment
X18079 N18079 N18080 Segment
X18080 N18080 N18081 Segment
X18081 N18081 N18082 Segment
X18082 N18082 N18083 Segment
X18083 N18083 N18084 Segment
X18084 N18084 N18085 Segment
X18085 N18085 N18086 Segment
X18086 N18086 N18087 Segment
X18087 N18087 N18088 Segment
X18088 N18088 N18089 Segment
X18089 N18089 N18090 Segment
X18090 N18090 N18091 Segment
X18091 N18091 N18092 Segment
X18092 N18092 N18093 Segment
X18093 N18093 N18094 Segment
X18094 N18094 N18095 Segment
X18095 N18095 N18096 Segment
X18096 N18096 N18097 Segment
X18097 N18097 N18098 Segment
X18098 N18098 N18099 Segment
X18099 N18099 N18100 Segment
X18100 N18100 N18101 Segment
X18101 N18101 N18102 Segment
X18102 N18102 N18103 Segment
X18103 N18103 N18104 Segment
X18104 N18104 N18105 Segment
X18105 N18105 N18106 Segment
X18106 N18106 N18107 Segment
X18107 N18107 N18108 Segment
X18108 N18108 N18109 Segment
X18109 N18109 N18110 Segment
X18110 N18110 N18111 Segment
X18111 N18111 N18112 Segment
X18112 N18112 N18113 Segment
X18113 N18113 N18114 Segment
X18114 N18114 N18115 Segment
X18115 N18115 N18116 Segment
X18116 N18116 N18117 Segment
X18117 N18117 N18118 Segment
X18118 N18118 N18119 Segment
X18119 N18119 N18120 Segment
X18120 N18120 N18121 Segment
X18121 N18121 N18122 Segment
X18122 N18122 N18123 Segment
X18123 N18123 N18124 Segment
X18124 N18124 N18125 Segment
X18125 N18125 N18126 Segment
X18126 N18126 N18127 Segment
X18127 N18127 N18128 Segment
X18128 N18128 N18129 Segment
X18129 N18129 N18130 Segment
X18130 N18130 N18131 Segment
X18131 N18131 N18132 Segment
X18132 N18132 N18133 Segment
X18133 N18133 N18134 Segment
X18134 N18134 N18135 Segment
X18135 N18135 N18136 Segment
X18136 N18136 N18137 Segment
X18137 N18137 N18138 Segment
X18138 N18138 N18139 Segment
X18139 N18139 N18140 Segment
X18140 N18140 N18141 Segment
X18141 N18141 N18142 Segment
X18142 N18142 N18143 Segment
X18143 N18143 N18144 Segment
X18144 N18144 N18145 Segment
X18145 N18145 N18146 Segment
X18146 N18146 N18147 Segment
X18147 N18147 N18148 Segment
X18148 N18148 N18149 Segment
X18149 N18149 N18150 Segment
X18150 N18150 N18151 Segment
X18151 N18151 N18152 Segment
X18152 N18152 N18153 Segment
X18153 N18153 N18154 Segment
X18154 N18154 N18155 Segment
X18155 N18155 N18156 Segment
X18156 N18156 N18157 Segment
X18157 N18157 N18158 Segment
X18158 N18158 N18159 Segment
X18159 N18159 N18160 Segment
X18160 N18160 N18161 Segment
X18161 N18161 N18162 Segment
X18162 N18162 N18163 Segment
X18163 N18163 N18164 Segment
X18164 N18164 N18165 Segment
X18165 N18165 N18166 Segment
X18166 N18166 N18167 Segment
X18167 N18167 N18168 Segment
X18168 N18168 N18169 Segment
X18169 N18169 N18170 Segment
X18170 N18170 N18171 Segment
X18171 N18171 N18172 Segment
X18172 N18172 N18173 Segment
X18173 N18173 N18174 Segment
X18174 N18174 N18175 Segment
X18175 N18175 N18176 Segment
X18176 N18176 N18177 Segment
X18177 N18177 N18178 Segment
X18178 N18178 N18179 Segment
X18179 N18179 N18180 Segment
X18180 N18180 N18181 Segment
X18181 N18181 N18182 Segment
X18182 N18182 N18183 Segment
X18183 N18183 N18184 Segment
X18184 N18184 N18185 Segment
X18185 N18185 N18186 Segment
X18186 N18186 N18187 Segment
X18187 N18187 N18188 Segment
X18188 N18188 N18189 Segment
X18189 N18189 N18190 Segment
X18190 N18190 N18191 Segment
X18191 N18191 N18192 Segment
X18192 N18192 N18193 Segment
X18193 N18193 N18194 Segment
X18194 N18194 N18195 Segment
X18195 N18195 N18196 Segment
X18196 N18196 N18197 Segment
X18197 N18197 N18198 Segment
X18198 N18198 N18199 Segment
X18199 N18199 N18200 Segment
X18200 N18200 N18201 Segment
X18201 N18201 N18202 Segment
X18202 N18202 N18203 Segment
X18203 N18203 N18204 Segment
X18204 N18204 N18205 Segment
X18205 N18205 N18206 Segment
X18206 N18206 N18207 Segment
X18207 N18207 N18208 Segment
X18208 N18208 N18209 Segment
X18209 N18209 N18210 Segment
X18210 N18210 N18211 Segment
X18211 N18211 N18212 Segment
X18212 N18212 N18213 Segment
X18213 N18213 N18214 Segment
X18214 N18214 N18215 Segment
X18215 N18215 N18216 Segment
X18216 N18216 N18217 Segment
X18217 N18217 N18218 Segment
X18218 N18218 N18219 Segment
X18219 N18219 N18220 Segment
X18220 N18220 N18221 Segment
X18221 N18221 N18222 Segment
X18222 N18222 N18223 Segment
X18223 N18223 N18224 Segment
X18224 N18224 N18225 Segment
X18225 N18225 N18226 Segment
X18226 N18226 N18227 Segment
X18227 N18227 N18228 Segment
X18228 N18228 N18229 Segment
X18229 N18229 N18230 Segment
X18230 N18230 N18231 Segment
X18231 N18231 N18232 Segment
X18232 N18232 N18233 Segment
X18233 N18233 N18234 Segment
X18234 N18234 N18235 Segment
X18235 N18235 N18236 Segment
X18236 N18236 N18237 Segment
X18237 N18237 N18238 Segment
X18238 N18238 N18239 Segment
X18239 N18239 N18240 Segment
X18240 N18240 N18241 Segment
X18241 N18241 N18242 Segment
X18242 N18242 N18243 Segment
X18243 N18243 N18244 Segment
X18244 N18244 N18245 Segment
X18245 N18245 N18246 Segment
X18246 N18246 N18247 Segment
X18247 N18247 N18248 Segment
X18248 N18248 N18249 Segment
X18249 N18249 N18250 Segment
X18250 N18250 N18251 Segment
X18251 N18251 N18252 Segment
X18252 N18252 N18253 Segment
X18253 N18253 N18254 Segment
X18254 N18254 N18255 Segment
X18255 N18255 N18256 Segment
X18256 N18256 N18257 Segment
X18257 N18257 N18258 Segment
X18258 N18258 N18259 Segment
X18259 N18259 N18260 Segment
X18260 N18260 N18261 Segment
X18261 N18261 N18262 Segment
X18262 N18262 N18263 Segment
X18263 N18263 N18264 Segment
X18264 N18264 N18265 Segment
X18265 N18265 N18266 Segment
X18266 N18266 N18267 Segment
X18267 N18267 N18268 Segment
X18268 N18268 N18269 Segment
X18269 N18269 N18270 Segment
X18270 N18270 N18271 Segment
X18271 N18271 N18272 Segment
X18272 N18272 N18273 Segment
X18273 N18273 N18274 Segment
X18274 N18274 N18275 Segment
X18275 N18275 N18276 Segment
X18276 N18276 N18277 Segment
X18277 N18277 N18278 Segment
X18278 N18278 N18279 Segment
X18279 N18279 N18280 Segment
X18280 N18280 N18281 Segment
X18281 N18281 N18282 Segment
X18282 N18282 N18283 Segment
X18283 N18283 N18284 Segment
X18284 N18284 N18285 Segment
X18285 N18285 N18286 Segment
X18286 N18286 N18287 Segment
X18287 N18287 N18288 Segment
X18288 N18288 N18289 Segment
X18289 N18289 N18290 Segment
X18290 N18290 N18291 Segment
X18291 N18291 N18292 Segment
X18292 N18292 N18293 Segment
X18293 N18293 N18294 Segment
X18294 N18294 N18295 Segment
X18295 N18295 N18296 Segment
X18296 N18296 N18297 Segment
X18297 N18297 N18298 Segment
X18298 N18298 N18299 Segment
X18299 N18299 N18300 Segment
X18300 N18300 N18301 Segment
X18301 N18301 N18302 Segment
X18302 N18302 N18303 Segment
X18303 N18303 N18304 Segment
X18304 N18304 N18305 Segment
X18305 N18305 N18306 Segment
X18306 N18306 N18307 Segment
X18307 N18307 N18308 Segment
X18308 N18308 N18309 Segment
X18309 N18309 N18310 Segment
X18310 N18310 N18311 Segment
X18311 N18311 N18312 Segment
X18312 N18312 N18313 Segment
X18313 N18313 N18314 Segment
X18314 N18314 N18315 Segment
X18315 N18315 N18316 Segment
X18316 N18316 N18317 Segment
X18317 N18317 N18318 Segment
X18318 N18318 N18319 Segment
X18319 N18319 N18320 Segment
X18320 N18320 N18321 Segment
X18321 N18321 N18322 Segment
X18322 N18322 N18323 Segment
X18323 N18323 N18324 Segment
X18324 N18324 N18325 Segment
X18325 N18325 N18326 Segment
X18326 N18326 N18327 Segment
X18327 N18327 N18328 Segment
X18328 N18328 N18329 Segment
X18329 N18329 N18330 Segment
X18330 N18330 N18331 Segment
X18331 N18331 N18332 Segment
X18332 N18332 N18333 Segment
X18333 N18333 N18334 Segment
X18334 N18334 N18335 Segment
X18335 N18335 N18336 Segment
X18336 N18336 N18337 Segment
X18337 N18337 N18338 Segment
X18338 N18338 N18339 Segment
X18339 N18339 N18340 Segment
X18340 N18340 N18341 Segment
X18341 N18341 N18342 Segment
X18342 N18342 N18343 Segment
X18343 N18343 N18344 Segment
X18344 N18344 N18345 Segment
X18345 N18345 N18346 Segment
X18346 N18346 N18347 Segment
X18347 N18347 N18348 Segment
X18348 N18348 N18349 Segment
X18349 N18349 N18350 Segment
X18350 N18350 N18351 Segment
X18351 N18351 N18352 Segment
X18352 N18352 N18353 Segment
X18353 N18353 N18354 Segment
X18354 N18354 N18355 Segment
X18355 N18355 N18356 Segment
X18356 N18356 N18357 Segment
X18357 N18357 N18358 Segment
X18358 N18358 N18359 Segment
X18359 N18359 N18360 Segment
X18360 N18360 N18361 Segment
X18361 N18361 N18362 Segment
X18362 N18362 N18363 Segment
X18363 N18363 N18364 Segment
X18364 N18364 N18365 Segment
X18365 N18365 N18366 Segment
X18366 N18366 N18367 Segment
X18367 N18367 N18368 Segment
X18368 N18368 N18369 Segment
X18369 N18369 N18370 Segment
X18370 N18370 N18371 Segment
X18371 N18371 N18372 Segment
X18372 N18372 N18373 Segment
X18373 N18373 N18374 Segment
X18374 N18374 N18375 Segment
X18375 N18375 N18376 Segment
X18376 N18376 N18377 Segment
X18377 N18377 N18378 Segment
X18378 N18378 N18379 Segment
X18379 N18379 N18380 Segment
X18380 N18380 N18381 Segment
X18381 N18381 N18382 Segment
X18382 N18382 N18383 Segment
X18383 N18383 N18384 Segment
X18384 N18384 N18385 Segment
X18385 N18385 N18386 Segment
X18386 N18386 N18387 Segment
X18387 N18387 N18388 Segment
X18388 N18388 N18389 Segment
X18389 N18389 N18390 Segment
X18390 N18390 N18391 Segment
X18391 N18391 N18392 Segment
X18392 N18392 N18393 Segment
X18393 N18393 N18394 Segment
X18394 N18394 N18395 Segment
X18395 N18395 N18396 Segment
X18396 N18396 N18397 Segment
X18397 N18397 N18398 Segment
X18398 N18398 N18399 Segment
X18399 N18399 N18400 Segment
X18400 N18400 N18401 Segment
X18401 N18401 N18402 Segment
X18402 N18402 N18403 Segment
X18403 N18403 N18404 Segment
X18404 N18404 N18405 Segment
X18405 N18405 N18406 Segment
X18406 N18406 N18407 Segment
X18407 N18407 N18408 Segment
X18408 N18408 N18409 Segment
X18409 N18409 N18410 Segment
X18410 N18410 N18411 Segment
X18411 N18411 N18412 Segment
X18412 N18412 N18413 Segment
X18413 N18413 N18414 Segment
X18414 N18414 N18415 Segment
X18415 N18415 N18416 Segment
X18416 N18416 N18417 Segment
X18417 N18417 N18418 Segment
X18418 N18418 N18419 Segment
X18419 N18419 N18420 Segment
X18420 N18420 N18421 Segment
X18421 N18421 N18422 Segment
X18422 N18422 N18423 Segment
X18423 N18423 N18424 Segment
X18424 N18424 N18425 Segment
X18425 N18425 N18426 Segment
X18426 N18426 N18427 Segment
X18427 N18427 N18428 Segment
X18428 N18428 N18429 Segment
X18429 N18429 N18430 Segment
X18430 N18430 N18431 Segment
X18431 N18431 N18432 Segment
X18432 N18432 N18433 Segment
X18433 N18433 N18434 Segment
X18434 N18434 N18435 Segment
X18435 N18435 N18436 Segment
X18436 N18436 N18437 Segment
X18437 N18437 N18438 Segment
X18438 N18438 N18439 Segment
X18439 N18439 N18440 Segment
X18440 N18440 N18441 Segment
X18441 N18441 N18442 Segment
X18442 N18442 N18443 Segment
X18443 N18443 N18444 Segment
X18444 N18444 N18445 Segment
X18445 N18445 N18446 Segment
X18446 N18446 N18447 Segment
X18447 N18447 N18448 Segment
X18448 N18448 N18449 Segment
X18449 N18449 N18450 Segment
X18450 N18450 N18451 Segment
X18451 N18451 N18452 Segment
X18452 N18452 N18453 Segment
X18453 N18453 N18454 Segment
X18454 N18454 N18455 Segment
X18455 N18455 N18456 Segment
X18456 N18456 N18457 Segment
X18457 N18457 N18458 Segment
X18458 N18458 N18459 Segment
X18459 N18459 N18460 Segment
X18460 N18460 N18461 Segment
X18461 N18461 N18462 Segment
X18462 N18462 N18463 Segment
X18463 N18463 N18464 Segment
X18464 N18464 N18465 Segment
X18465 N18465 N18466 Segment
X18466 N18466 N18467 Segment
X18467 N18467 N18468 Segment
X18468 N18468 N18469 Segment
X18469 N18469 N18470 Segment
X18470 N18470 N18471 Segment
X18471 N18471 N18472 Segment
X18472 N18472 N18473 Segment
X18473 N18473 N18474 Segment
X18474 N18474 N18475 Segment
X18475 N18475 N18476 Segment
X18476 N18476 N18477 Segment
X18477 N18477 N18478 Segment
X18478 N18478 N18479 Segment
X18479 N18479 N18480 Segment
X18480 N18480 N18481 Segment
X18481 N18481 N18482 Segment
X18482 N18482 N18483 Segment
X18483 N18483 N18484 Segment
X18484 N18484 N18485 Segment
X18485 N18485 N18486 Segment
X18486 N18486 N18487 Segment
X18487 N18487 N18488 Segment
X18488 N18488 N18489 Segment
X18489 N18489 N18490 Segment
X18490 N18490 N18491 Segment
X18491 N18491 N18492 Segment
X18492 N18492 N18493 Segment
X18493 N18493 N18494 Segment
X18494 N18494 N18495 Segment
X18495 N18495 N18496 Segment
X18496 N18496 N18497 Segment
X18497 N18497 N18498 Segment
X18498 N18498 N18499 Segment
X18499 N18499 N18500 Segment
X18500 N18500 N18501 Segment
X18501 N18501 N18502 Segment
X18502 N18502 N18503 Segment
X18503 N18503 N18504 Segment
X18504 N18504 N18505 Segment
X18505 N18505 N18506 Segment
X18506 N18506 N18507 Segment
X18507 N18507 N18508 Segment
X18508 N18508 N18509 Segment
X18509 N18509 N18510 Segment
X18510 N18510 N18511 Segment
X18511 N18511 N18512 Segment
X18512 N18512 N18513 Segment
X18513 N18513 N18514 Segment
X18514 N18514 N18515 Segment
X18515 N18515 N18516 Segment
X18516 N18516 N18517 Segment
X18517 N18517 N18518 Segment
X18518 N18518 N18519 Segment
X18519 N18519 N18520 Segment
X18520 N18520 N18521 Segment
X18521 N18521 N18522 Segment
X18522 N18522 N18523 Segment
X18523 N18523 N18524 Segment
X18524 N18524 N18525 Segment
X18525 N18525 N18526 Segment
X18526 N18526 N18527 Segment
X18527 N18527 N18528 Segment
X18528 N18528 N18529 Segment
X18529 N18529 N18530 Segment
X18530 N18530 N18531 Segment
X18531 N18531 N18532 Segment
X18532 N18532 N18533 Segment
X18533 N18533 N18534 Segment
X18534 N18534 N18535 Segment
X18535 N18535 N18536 Segment
X18536 N18536 N18537 Segment
X18537 N18537 N18538 Segment
X18538 N18538 N18539 Segment
X18539 N18539 N18540 Segment
X18540 N18540 N18541 Segment
X18541 N18541 N18542 Segment
X18542 N18542 N18543 Segment
X18543 N18543 N18544 Segment
X18544 N18544 N18545 Segment
X18545 N18545 N18546 Segment
X18546 N18546 N18547 Segment
X18547 N18547 N18548 Segment
X18548 N18548 N18549 Segment
X18549 N18549 N18550 Segment
X18550 N18550 N18551 Segment
X18551 N18551 N18552 Segment
X18552 N18552 N18553 Segment
X18553 N18553 N18554 Segment
X18554 N18554 N18555 Segment
X18555 N18555 N18556 Segment
X18556 N18556 N18557 Segment
X18557 N18557 N18558 Segment
X18558 N18558 N18559 Segment
X18559 N18559 N18560 Segment
X18560 N18560 N18561 Segment
X18561 N18561 N18562 Segment
X18562 N18562 N18563 Segment
X18563 N18563 N18564 Segment
X18564 N18564 N18565 Segment
X18565 N18565 N18566 Segment
X18566 N18566 N18567 Segment
X18567 N18567 N18568 Segment
X18568 N18568 N18569 Segment
X18569 N18569 N18570 Segment
X18570 N18570 N18571 Segment
X18571 N18571 N18572 Segment
X18572 N18572 N18573 Segment
X18573 N18573 N18574 Segment
X18574 N18574 N18575 Segment
X18575 N18575 N18576 Segment
X18576 N18576 N18577 Segment
X18577 N18577 N18578 Segment
X18578 N18578 N18579 Segment
X18579 N18579 N18580 Segment
X18580 N18580 N18581 Segment
X18581 N18581 N18582 Segment
X18582 N18582 N18583 Segment
X18583 N18583 N18584 Segment
X18584 N18584 N18585 Segment
X18585 N18585 N18586 Segment
X18586 N18586 N18587 Segment
X18587 N18587 N18588 Segment
X18588 N18588 N18589 Segment
X18589 N18589 N18590 Segment
X18590 N18590 N18591 Segment
X18591 N18591 N18592 Segment
X18592 N18592 N18593 Segment
X18593 N18593 N18594 Segment
X18594 N18594 N18595 Segment
X18595 N18595 N18596 Segment
X18596 N18596 N18597 Segment
X18597 N18597 N18598 Segment
X18598 N18598 N18599 Segment
X18599 N18599 N18600 Segment
X18600 N18600 N18601 Segment
X18601 N18601 N18602 Segment
X18602 N18602 N18603 Segment
X18603 N18603 N18604 Segment
X18604 N18604 N18605 Segment
X18605 N18605 N18606 Segment
X18606 N18606 N18607 Segment
X18607 N18607 N18608 Segment
X18608 N18608 N18609 Segment
X18609 N18609 N18610 Segment
X18610 N18610 N18611 Segment
X18611 N18611 N18612 Segment
X18612 N18612 N18613 Segment
X18613 N18613 N18614 Segment
X18614 N18614 N18615 Segment
X18615 N18615 N18616 Segment
X18616 N18616 N18617 Segment
X18617 N18617 N18618 Segment
X18618 N18618 N18619 Segment
X18619 N18619 N18620 Segment
X18620 N18620 N18621 Segment
X18621 N18621 N18622 Segment
X18622 N18622 N18623 Segment
X18623 N18623 N18624 Segment
X18624 N18624 N18625 Segment
X18625 N18625 N18626 Segment
X18626 N18626 N18627 Segment
X18627 N18627 N18628 Segment
X18628 N18628 N18629 Segment
X18629 N18629 N18630 Segment
X18630 N18630 N18631 Segment
X18631 N18631 N18632 Segment
X18632 N18632 N18633 Segment
X18633 N18633 N18634 Segment
X18634 N18634 N18635 Segment
X18635 N18635 N18636 Segment
X18636 N18636 N18637 Segment
X18637 N18637 N18638 Segment
X18638 N18638 N18639 Segment
X18639 N18639 N18640 Segment
X18640 N18640 N18641 Segment
X18641 N18641 N18642 Segment
X18642 N18642 N18643 Segment
X18643 N18643 N18644 Segment
X18644 N18644 N18645 Segment
X18645 N18645 N18646 Segment
X18646 N18646 N18647 Segment
X18647 N18647 N18648 Segment
X18648 N18648 N18649 Segment
X18649 N18649 N18650 Segment
X18650 N18650 N18651 Segment
X18651 N18651 N18652 Segment
X18652 N18652 N18653 Segment
X18653 N18653 N18654 Segment
X18654 N18654 N18655 Segment
X18655 N18655 N18656 Segment
X18656 N18656 N18657 Segment
X18657 N18657 N18658 Segment
X18658 N18658 N18659 Segment
X18659 N18659 N18660 Segment
X18660 N18660 N18661 Segment
X18661 N18661 N18662 Segment
X18662 N18662 N18663 Segment
X18663 N18663 N18664 Segment
X18664 N18664 N18665 Segment
X18665 N18665 N18666 Segment
X18666 N18666 N18667 Segment
X18667 N18667 N18668 Segment
X18668 N18668 N18669 Segment
X18669 N18669 N18670 Segment
X18670 N18670 N18671 Segment
X18671 N18671 N18672 Segment
X18672 N18672 N18673 Segment
X18673 N18673 N18674 Segment
X18674 N18674 N18675 Segment
X18675 N18675 N18676 Segment
X18676 N18676 N18677 Segment
X18677 N18677 N18678 Segment
X18678 N18678 N18679 Segment
X18679 N18679 N18680 Segment
X18680 N18680 N18681 Segment
X18681 N18681 N18682 Segment
X18682 N18682 N18683 Segment
X18683 N18683 N18684 Segment
X18684 N18684 N18685 Segment
X18685 N18685 N18686 Segment
X18686 N18686 N18687 Segment
X18687 N18687 N18688 Segment
X18688 N18688 N18689 Segment
X18689 N18689 N18690 Segment
X18690 N18690 N18691 Segment
X18691 N18691 N18692 Segment
X18692 N18692 N18693 Segment
X18693 N18693 N18694 Segment
X18694 N18694 N18695 Segment
X18695 N18695 N18696 Segment
X18696 N18696 N18697 Segment
X18697 N18697 N18698 Segment
X18698 N18698 N18699 Segment
X18699 N18699 N18700 Segment
X18700 N18700 N18701 Segment
X18701 N18701 N18702 Segment
X18702 N18702 N18703 Segment
X18703 N18703 N18704 Segment
X18704 N18704 N18705 Segment
X18705 N18705 N18706 Segment
X18706 N18706 N18707 Segment
X18707 N18707 N18708 Segment
X18708 N18708 N18709 Segment
X18709 N18709 N18710 Segment
X18710 N18710 N18711 Segment
X18711 N18711 N18712 Segment
X18712 N18712 N18713 Segment
X18713 N18713 N18714 Segment
X18714 N18714 N18715 Segment
X18715 N18715 N18716 Segment
X18716 N18716 N18717 Segment
X18717 N18717 N18718 Segment
X18718 N18718 N18719 Segment
X18719 N18719 N18720 Segment
X18720 N18720 N18721 Segment
X18721 N18721 N18722 Segment
X18722 N18722 N18723 Segment
X18723 N18723 N18724 Segment
X18724 N18724 N18725 Segment
X18725 N18725 N18726 Segment
X18726 N18726 N18727 Segment
X18727 N18727 N18728 Segment
X18728 N18728 N18729 Segment
X18729 N18729 N18730 Segment
X18730 N18730 N18731 Segment
X18731 N18731 N18732 Segment
X18732 N18732 N18733 Segment
X18733 N18733 N18734 Segment
X18734 N18734 N18735 Segment
X18735 N18735 N18736 Segment
X18736 N18736 N18737 Segment
X18737 N18737 N18738 Segment
X18738 N18738 N18739 Segment
X18739 N18739 N18740 Segment
X18740 N18740 N18741 Segment
X18741 N18741 N18742 Segment
X18742 N18742 N18743 Segment
X18743 N18743 N18744 Segment
X18744 N18744 N18745 Segment
X18745 N18745 N18746 Segment
X18746 N18746 N18747 Segment
X18747 N18747 N18748 Segment
X18748 N18748 N18749 Segment
X18749 N18749 N18750 Segment
X18750 N18750 N18751 Segment
X18751 N18751 N18752 Segment
X18752 N18752 N18753 Segment
X18753 N18753 N18754 Segment
X18754 N18754 N18755 Segment
X18755 N18755 N18756 Segment
X18756 N18756 N18757 Segment
X18757 N18757 N18758 Segment
X18758 N18758 N18759 Segment
X18759 N18759 N18760 Segment
X18760 N18760 N18761 Segment
X18761 N18761 N18762 Segment
X18762 N18762 N18763 Segment
X18763 N18763 N18764 Segment
X18764 N18764 N18765 Segment
X18765 N18765 N18766 Segment
X18766 N18766 N18767 Segment
X18767 N18767 N18768 Segment
X18768 N18768 N18769 Segment
X18769 N18769 N18770 Segment
X18770 N18770 N18771 Segment
X18771 N18771 N18772 Segment
X18772 N18772 N18773 Segment
X18773 N18773 N18774 Segment
X18774 N18774 N18775 Segment
X18775 N18775 N18776 Segment
X18776 N18776 N18777 Segment
X18777 N18777 N18778 Segment
X18778 N18778 N18779 Segment
X18779 N18779 N18780 Segment
X18780 N18780 N18781 Segment
X18781 N18781 N18782 Segment
X18782 N18782 N18783 Segment
X18783 N18783 N18784 Segment
X18784 N18784 N18785 Segment
X18785 N18785 N18786 Segment
X18786 N18786 N18787 Segment
X18787 N18787 N18788 Segment
X18788 N18788 N18789 Segment
X18789 N18789 N18790 Segment
X18790 N18790 N18791 Segment
X18791 N18791 N18792 Segment
X18792 N18792 N18793 Segment
X18793 N18793 N18794 Segment
X18794 N18794 N18795 Segment
X18795 N18795 N18796 Segment
X18796 N18796 N18797 Segment
X18797 N18797 N18798 Segment
X18798 N18798 N18799 Segment
X18799 N18799 N18800 Segment
X18800 N18800 N18801 Segment
X18801 N18801 N18802 Segment
X18802 N18802 N18803 Segment
X18803 N18803 N18804 Segment
X18804 N18804 N18805 Segment
X18805 N18805 N18806 Segment
X18806 N18806 N18807 Segment
X18807 N18807 N18808 Segment
X18808 N18808 N18809 Segment
X18809 N18809 N18810 Segment
X18810 N18810 N18811 Segment
X18811 N18811 N18812 Segment
X18812 N18812 N18813 Segment
X18813 N18813 N18814 Segment
X18814 N18814 N18815 Segment
X18815 N18815 N18816 Segment
X18816 N18816 N18817 Segment
X18817 N18817 N18818 Segment
X18818 N18818 N18819 Segment
X18819 N18819 N18820 Segment
X18820 N18820 N18821 Segment
X18821 N18821 N18822 Segment
X18822 N18822 N18823 Segment
X18823 N18823 N18824 Segment
X18824 N18824 N18825 Segment
X18825 N18825 N18826 Segment
X18826 N18826 N18827 Segment
X18827 N18827 N18828 Segment
X18828 N18828 N18829 Segment
X18829 N18829 N18830 Segment
X18830 N18830 N18831 Segment
X18831 N18831 N18832 Segment
X18832 N18832 N18833 Segment
X18833 N18833 N18834 Segment
X18834 N18834 N18835 Segment
X18835 N18835 N18836 Segment
X18836 N18836 N18837 Segment
X18837 N18837 N18838 Segment
X18838 N18838 N18839 Segment
X18839 N18839 N18840 Segment
X18840 N18840 N18841 Segment
X18841 N18841 N18842 Segment
X18842 N18842 N18843 Segment
X18843 N18843 N18844 Segment
X18844 N18844 N18845 Segment
X18845 N18845 N18846 Segment
X18846 N18846 N18847 Segment
X18847 N18847 N18848 Segment
X18848 N18848 N18849 Segment
X18849 N18849 N18850 Segment
X18850 N18850 N18851 Segment
X18851 N18851 N18852 Segment
X18852 N18852 N18853 Segment
X18853 N18853 N18854 Segment
X18854 N18854 N18855 Segment
X18855 N18855 N18856 Segment
X18856 N18856 N18857 Segment
X18857 N18857 N18858 Segment
X18858 N18858 N18859 Segment
X18859 N18859 N18860 Segment
X18860 N18860 N18861 Segment
X18861 N18861 N18862 Segment
X18862 N18862 N18863 Segment
X18863 N18863 N18864 Segment
X18864 N18864 N18865 Segment
X18865 N18865 N18866 Segment
X18866 N18866 N18867 Segment
X18867 N18867 N18868 Segment
X18868 N18868 N18869 Segment
X18869 N18869 N18870 Segment
X18870 N18870 N18871 Segment
X18871 N18871 N18872 Segment
X18872 N18872 N18873 Segment
X18873 N18873 N18874 Segment
X18874 N18874 N18875 Segment
X18875 N18875 N18876 Segment
X18876 N18876 N18877 Segment
X18877 N18877 N18878 Segment
X18878 N18878 N18879 Segment
X18879 N18879 N18880 Segment
X18880 N18880 N18881 Segment
X18881 N18881 N18882 Segment
X18882 N18882 N18883 Segment
X18883 N18883 N18884 Segment
X18884 N18884 N18885 Segment
X18885 N18885 N18886 Segment
X18886 N18886 N18887 Segment
X18887 N18887 N18888 Segment
X18888 N18888 N18889 Segment
X18889 N18889 N18890 Segment
X18890 N18890 N18891 Segment
X18891 N18891 N18892 Segment
X18892 N18892 N18893 Segment
X18893 N18893 N18894 Segment
X18894 N18894 N18895 Segment
X18895 N18895 N18896 Segment
X18896 N18896 N18897 Segment
X18897 N18897 N18898 Segment
X18898 N18898 N18899 Segment
X18899 N18899 N18900 Segment
X18900 N18900 N18901 Segment
X18901 N18901 N18902 Segment
X18902 N18902 N18903 Segment
X18903 N18903 N18904 Segment
X18904 N18904 N18905 Segment
X18905 N18905 N18906 Segment
X18906 N18906 N18907 Segment
X18907 N18907 N18908 Segment
X18908 N18908 N18909 Segment
X18909 N18909 N18910 Segment
X18910 N18910 N18911 Segment
X18911 N18911 N18912 Segment
X18912 N18912 N18913 Segment
X18913 N18913 N18914 Segment
X18914 N18914 N18915 Segment
X18915 N18915 N18916 Segment
X18916 N18916 N18917 Segment
X18917 N18917 N18918 Segment
X18918 N18918 N18919 Segment
X18919 N18919 N18920 Segment
X18920 N18920 N18921 Segment
X18921 N18921 N18922 Segment
X18922 N18922 N18923 Segment
X18923 N18923 N18924 Segment
X18924 N18924 N18925 Segment
X18925 N18925 N18926 Segment
X18926 N18926 N18927 Segment
X18927 N18927 N18928 Segment
X18928 N18928 N18929 Segment
X18929 N18929 N18930 Segment
X18930 N18930 N18931 Segment
X18931 N18931 N18932 Segment
X18932 N18932 N18933 Segment
X18933 N18933 N18934 Segment
X18934 N18934 N18935 Segment
X18935 N18935 N18936 Segment
X18936 N18936 N18937 Segment
X18937 N18937 N18938 Segment
X18938 N18938 N18939 Segment
X18939 N18939 N18940 Segment
X18940 N18940 N18941 Segment
X18941 N18941 N18942 Segment
X18942 N18942 N18943 Segment
X18943 N18943 N18944 Segment
X18944 N18944 N18945 Segment
X18945 N18945 N18946 Segment
X18946 N18946 N18947 Segment
X18947 N18947 N18948 Segment
X18948 N18948 N18949 Segment
X18949 N18949 N18950 Segment
X18950 N18950 N18951 Segment
X18951 N18951 N18952 Segment
X18952 N18952 N18953 Segment
X18953 N18953 N18954 Segment
X18954 N18954 N18955 Segment
X18955 N18955 N18956 Segment
X18956 N18956 N18957 Segment
X18957 N18957 N18958 Segment
X18958 N18958 N18959 Segment
X18959 N18959 N18960 Segment
X18960 N18960 N18961 Segment
X18961 N18961 N18962 Segment
X18962 N18962 N18963 Segment
X18963 N18963 N18964 Segment
X18964 N18964 N18965 Segment
X18965 N18965 N18966 Segment
X18966 N18966 N18967 Segment
X18967 N18967 N18968 Segment
X18968 N18968 N18969 Segment
X18969 N18969 N18970 Segment
X18970 N18970 N18971 Segment
X18971 N18971 N18972 Segment
X18972 N18972 N18973 Segment
X18973 N18973 N18974 Segment
X18974 N18974 N18975 Segment
X18975 N18975 N18976 Segment
X18976 N18976 N18977 Segment
X18977 N18977 N18978 Segment
X18978 N18978 N18979 Segment
X18979 N18979 N18980 Segment
X18980 N18980 N18981 Segment
X18981 N18981 N18982 Segment
X18982 N18982 N18983 Segment
X18983 N18983 N18984 Segment
X18984 N18984 N18985 Segment
X18985 N18985 N18986 Segment
X18986 N18986 N18987 Segment
X18987 N18987 N18988 Segment
X18988 N18988 N18989 Segment
X18989 N18989 N18990 Segment
X18990 N18990 N18991 Segment
X18991 N18991 N18992 Segment
X18992 N18992 N18993 Segment
X18993 N18993 N18994 Segment
X18994 N18994 N18995 Segment
X18995 N18995 N18996 Segment
X18996 N18996 N18997 Segment
X18997 N18997 N18998 Segment
X18998 N18998 N18999 Segment
X18999 N18999 N19000 Segment
X19000 N19000 N19001 Segment
X19001 N19001 N19002 Segment
X19002 N19002 N19003 Segment
X19003 N19003 N19004 Segment
X19004 N19004 N19005 Segment
X19005 N19005 N19006 Segment
X19006 N19006 N19007 Segment
X19007 N19007 N19008 Segment
X19008 N19008 N19009 Segment
X19009 N19009 N19010 Segment
X19010 N19010 N19011 Segment
X19011 N19011 N19012 Segment
X19012 N19012 N19013 Segment
X19013 N19013 N19014 Segment
X19014 N19014 N19015 Segment
X19015 N19015 N19016 Segment
X19016 N19016 N19017 Segment
X19017 N19017 N19018 Segment
X19018 N19018 N19019 Segment
X19019 N19019 N19020 Segment
X19020 N19020 N19021 Segment
X19021 N19021 N19022 Segment
X19022 N19022 N19023 Segment
X19023 N19023 N19024 Segment
X19024 N19024 N19025 Segment
X19025 N19025 N19026 Segment
X19026 N19026 N19027 Segment
X19027 N19027 N19028 Segment
X19028 N19028 N19029 Segment
X19029 N19029 N19030 Segment
X19030 N19030 N19031 Segment
X19031 N19031 N19032 Segment
X19032 N19032 N19033 Segment
X19033 N19033 N19034 Segment
X19034 N19034 N19035 Segment
X19035 N19035 N19036 Segment
X19036 N19036 N19037 Segment
X19037 N19037 N19038 Segment
X19038 N19038 N19039 Segment
X19039 N19039 N19040 Segment
X19040 N19040 N19041 Segment
X19041 N19041 N19042 Segment
X19042 N19042 N19043 Segment
X19043 N19043 N19044 Segment
X19044 N19044 N19045 Segment
X19045 N19045 N19046 Segment
X19046 N19046 N19047 Segment
X19047 N19047 N19048 Segment
X19048 N19048 N19049 Segment
X19049 N19049 N19050 Segment
X19050 N19050 N19051 Segment
X19051 N19051 N19052 Segment
X19052 N19052 N19053 Segment
X19053 N19053 N19054 Segment
X19054 N19054 N19055 Segment
X19055 N19055 N19056 Segment
X19056 N19056 N19057 Segment
X19057 N19057 N19058 Segment
X19058 N19058 N19059 Segment
X19059 N19059 N19060 Segment
X19060 N19060 N19061 Segment
X19061 N19061 N19062 Segment
X19062 N19062 N19063 Segment
X19063 N19063 N19064 Segment
X19064 N19064 N19065 Segment
X19065 N19065 N19066 Segment
X19066 N19066 N19067 Segment
X19067 N19067 N19068 Segment
X19068 N19068 N19069 Segment
X19069 N19069 N19070 Segment
X19070 N19070 N19071 Segment
X19071 N19071 N19072 Segment
X19072 N19072 N19073 Segment
X19073 N19073 N19074 Segment
X19074 N19074 N19075 Segment
X19075 N19075 N19076 Segment
X19076 N19076 N19077 Segment
X19077 N19077 N19078 Segment
X19078 N19078 N19079 Segment
X19079 N19079 N19080 Segment
X19080 N19080 N19081 Segment
X19081 N19081 N19082 Segment
X19082 N19082 N19083 Segment
X19083 N19083 N19084 Segment
X19084 N19084 N19085 Segment
X19085 N19085 N19086 Segment
X19086 N19086 N19087 Segment
X19087 N19087 N19088 Segment
X19088 N19088 N19089 Segment
X19089 N19089 N19090 Segment
X19090 N19090 N19091 Segment
X19091 N19091 N19092 Segment
X19092 N19092 N19093 Segment
X19093 N19093 N19094 Segment
X19094 N19094 N19095 Segment
X19095 N19095 N19096 Segment
X19096 N19096 N19097 Segment
X19097 N19097 N19098 Segment
X19098 N19098 N19099 Segment
X19099 N19099 N19100 Segment
X19100 N19100 N19101 Segment
X19101 N19101 N19102 Segment
X19102 N19102 N19103 Segment
X19103 N19103 N19104 Segment
X19104 N19104 N19105 Segment
X19105 N19105 N19106 Segment
X19106 N19106 N19107 Segment
X19107 N19107 N19108 Segment
X19108 N19108 N19109 Segment
X19109 N19109 N19110 Segment
X19110 N19110 N19111 Segment
X19111 N19111 N19112 Segment
X19112 N19112 N19113 Segment
X19113 N19113 N19114 Segment
X19114 N19114 N19115 Segment
X19115 N19115 N19116 Segment
X19116 N19116 N19117 Segment
X19117 N19117 N19118 Segment
X19118 N19118 N19119 Segment
X19119 N19119 N19120 Segment
X19120 N19120 N19121 Segment
X19121 N19121 N19122 Segment
X19122 N19122 N19123 Segment
X19123 N19123 N19124 Segment
X19124 N19124 N19125 Segment
X19125 N19125 N19126 Segment
X19126 N19126 N19127 Segment
X19127 N19127 N19128 Segment
X19128 N19128 N19129 Segment
X19129 N19129 N19130 Segment
X19130 N19130 N19131 Segment
X19131 N19131 N19132 Segment
X19132 N19132 N19133 Segment
X19133 N19133 N19134 Segment
X19134 N19134 N19135 Segment
X19135 N19135 N19136 Segment
X19136 N19136 N19137 Segment
X19137 N19137 N19138 Segment
X19138 N19138 N19139 Segment
X19139 N19139 N19140 Segment
X19140 N19140 N19141 Segment
X19141 N19141 N19142 Segment
X19142 N19142 N19143 Segment
X19143 N19143 N19144 Segment
X19144 N19144 N19145 Segment
X19145 N19145 N19146 Segment
X19146 N19146 N19147 Segment
X19147 N19147 N19148 Segment
X19148 N19148 N19149 Segment
X19149 N19149 N19150 Segment
X19150 N19150 N19151 Segment
X19151 N19151 N19152 Segment
X19152 N19152 N19153 Segment
X19153 N19153 N19154 Segment
X19154 N19154 N19155 Segment
X19155 N19155 N19156 Segment
X19156 N19156 N19157 Segment
X19157 N19157 N19158 Segment
X19158 N19158 N19159 Segment
X19159 N19159 N19160 Segment
X19160 N19160 N19161 Segment
X19161 N19161 N19162 Segment
X19162 N19162 N19163 Segment
X19163 N19163 N19164 Segment
X19164 N19164 N19165 Segment
X19165 N19165 N19166 Segment
X19166 N19166 N19167 Segment
X19167 N19167 N19168 Segment
X19168 N19168 N19169 Segment
X19169 N19169 N19170 Segment
X19170 N19170 N19171 Segment
X19171 N19171 N19172 Segment
X19172 N19172 N19173 Segment
X19173 N19173 N19174 Segment
X19174 N19174 N19175 Segment
X19175 N19175 N19176 Segment
X19176 N19176 N19177 Segment
X19177 N19177 N19178 Segment
X19178 N19178 N19179 Segment
X19179 N19179 N19180 Segment
X19180 N19180 N19181 Segment
X19181 N19181 N19182 Segment
X19182 N19182 N19183 Segment
X19183 N19183 N19184 Segment
X19184 N19184 N19185 Segment
X19185 N19185 N19186 Segment
X19186 N19186 N19187 Segment
X19187 N19187 N19188 Segment
X19188 N19188 N19189 Segment
X19189 N19189 N19190 Segment
X19190 N19190 N19191 Segment
X19191 N19191 N19192 Segment
X19192 N19192 N19193 Segment
X19193 N19193 N19194 Segment
X19194 N19194 N19195 Segment
X19195 N19195 N19196 Segment
X19196 N19196 N19197 Segment
X19197 N19197 N19198 Segment
X19198 N19198 N19199 Segment
X19199 N19199 N19200 Segment
X19200 N19200 N19201 Segment
X19201 N19201 N19202 Segment
X19202 N19202 N19203 Segment
X19203 N19203 N19204 Segment
X19204 N19204 N19205 Segment
X19205 N19205 N19206 Segment
X19206 N19206 N19207 Segment
X19207 N19207 N19208 Segment
X19208 N19208 N19209 Segment
X19209 N19209 N19210 Segment
X19210 N19210 N19211 Segment
X19211 N19211 N19212 Segment
X19212 N19212 N19213 Segment
X19213 N19213 N19214 Segment
X19214 N19214 N19215 Segment
X19215 N19215 N19216 Segment
X19216 N19216 N19217 Segment
X19217 N19217 N19218 Segment
X19218 N19218 N19219 Segment
X19219 N19219 N19220 Segment
X19220 N19220 N19221 Segment
X19221 N19221 N19222 Segment
X19222 N19222 N19223 Segment
X19223 N19223 N19224 Segment
X19224 N19224 N19225 Segment
X19225 N19225 N19226 Segment
X19226 N19226 N19227 Segment
X19227 N19227 N19228 Segment
X19228 N19228 N19229 Segment
X19229 N19229 N19230 Segment
X19230 N19230 N19231 Segment
X19231 N19231 N19232 Segment
X19232 N19232 N19233 Segment
X19233 N19233 N19234 Segment
X19234 N19234 N19235 Segment
X19235 N19235 N19236 Segment
X19236 N19236 N19237 Segment
X19237 N19237 N19238 Segment
X19238 N19238 N19239 Segment
X19239 N19239 N19240 Segment
X19240 N19240 N19241 Segment
X19241 N19241 N19242 Segment
X19242 N19242 N19243 Segment
X19243 N19243 N19244 Segment
X19244 N19244 N19245 Segment
X19245 N19245 N19246 Segment
X19246 N19246 N19247 Segment
X19247 N19247 N19248 Segment
X19248 N19248 N19249 Segment
X19249 N19249 N19250 Segment
X19250 N19250 N19251 Segment
X19251 N19251 N19252 Segment
X19252 N19252 N19253 Segment
X19253 N19253 N19254 Segment
X19254 N19254 N19255 Segment
X19255 N19255 N19256 Segment
X19256 N19256 N19257 Segment
X19257 N19257 N19258 Segment
X19258 N19258 N19259 Segment
X19259 N19259 N19260 Segment
X19260 N19260 N19261 Segment
X19261 N19261 N19262 Segment
X19262 N19262 N19263 Segment
X19263 N19263 N19264 Segment
X19264 N19264 N19265 Segment
X19265 N19265 N19266 Segment
X19266 N19266 N19267 Segment
X19267 N19267 N19268 Segment
X19268 N19268 N19269 Segment
X19269 N19269 N19270 Segment
X19270 N19270 N19271 Segment
X19271 N19271 N19272 Segment
X19272 N19272 N19273 Segment
X19273 N19273 N19274 Segment
X19274 N19274 N19275 Segment
X19275 N19275 N19276 Segment
X19276 N19276 N19277 Segment
X19277 N19277 N19278 Segment
X19278 N19278 N19279 Segment
X19279 N19279 N19280 Segment
X19280 N19280 N19281 Segment
X19281 N19281 N19282 Segment
X19282 N19282 N19283 Segment
X19283 N19283 N19284 Segment
X19284 N19284 N19285 Segment
X19285 N19285 N19286 Segment
X19286 N19286 N19287 Segment
X19287 N19287 N19288 Segment
X19288 N19288 N19289 Segment
X19289 N19289 N19290 Segment
X19290 N19290 N19291 Segment
X19291 N19291 N19292 Segment
X19292 N19292 N19293 Segment
X19293 N19293 N19294 Segment
X19294 N19294 N19295 Segment
X19295 N19295 N19296 Segment
X19296 N19296 N19297 Segment
X19297 N19297 N19298 Segment
X19298 N19298 N19299 Segment
X19299 N19299 N19300 Segment
X19300 N19300 N19301 Segment
X19301 N19301 N19302 Segment
X19302 N19302 N19303 Segment
X19303 N19303 N19304 Segment
X19304 N19304 N19305 Segment
X19305 N19305 N19306 Segment
X19306 N19306 N19307 Segment
X19307 N19307 N19308 Segment
X19308 N19308 N19309 Segment
X19309 N19309 N19310 Segment
X19310 N19310 N19311 Segment
X19311 N19311 N19312 Segment
X19312 N19312 N19313 Segment
X19313 N19313 N19314 Segment
X19314 N19314 N19315 Segment
X19315 N19315 N19316 Segment
X19316 N19316 N19317 Segment
X19317 N19317 N19318 Segment
X19318 N19318 N19319 Segment
X19319 N19319 N19320 Segment
X19320 N19320 N19321 Segment
X19321 N19321 N19322 Segment
X19322 N19322 N19323 Segment
X19323 N19323 N19324 Segment
X19324 N19324 N19325 Segment
X19325 N19325 N19326 Segment
X19326 N19326 N19327 Segment
X19327 N19327 N19328 Segment
X19328 N19328 N19329 Segment
X19329 N19329 N19330 Segment
X19330 N19330 N19331 Segment
X19331 N19331 N19332 Segment
X19332 N19332 N19333 Segment
X19333 N19333 N19334 Segment
X19334 N19334 N19335 Segment
X19335 N19335 N19336 Segment
X19336 N19336 N19337 Segment
X19337 N19337 N19338 Segment
X19338 N19338 N19339 Segment
X19339 N19339 N19340 Segment
X19340 N19340 N19341 Segment
X19341 N19341 N19342 Segment
X19342 N19342 N19343 Segment
X19343 N19343 N19344 Segment
X19344 N19344 N19345 Segment
X19345 N19345 N19346 Segment
X19346 N19346 N19347 Segment
X19347 N19347 N19348 Segment
X19348 N19348 N19349 Segment
X19349 N19349 N19350 Segment
X19350 N19350 N19351 Segment
X19351 N19351 N19352 Segment
X19352 N19352 N19353 Segment
X19353 N19353 N19354 Segment
X19354 N19354 N19355 Segment
X19355 N19355 N19356 Segment
X19356 N19356 N19357 Segment
X19357 N19357 N19358 Segment
X19358 N19358 N19359 Segment
X19359 N19359 N19360 Segment
X19360 N19360 N19361 Segment
X19361 N19361 N19362 Segment
X19362 N19362 N19363 Segment
X19363 N19363 N19364 Segment
X19364 N19364 N19365 Segment
X19365 N19365 N19366 Segment
X19366 N19366 N19367 Segment
X19367 N19367 N19368 Segment
X19368 N19368 N19369 Segment
X19369 N19369 N19370 Segment
X19370 N19370 N19371 Segment
X19371 N19371 N19372 Segment
X19372 N19372 N19373 Segment
X19373 N19373 N19374 Segment
X19374 N19374 N19375 Segment
X19375 N19375 N19376 Segment
X19376 N19376 N19377 Segment
X19377 N19377 N19378 Segment
X19378 N19378 N19379 Segment
X19379 N19379 N19380 Segment
X19380 N19380 N19381 Segment
X19381 N19381 N19382 Segment
X19382 N19382 N19383 Segment
X19383 N19383 N19384 Segment
X19384 N19384 N19385 Segment
X19385 N19385 N19386 Segment
X19386 N19386 N19387 Segment
X19387 N19387 N19388 Segment
X19388 N19388 N19389 Segment
X19389 N19389 N19390 Segment
X19390 N19390 N19391 Segment
X19391 N19391 N19392 Segment
X19392 N19392 N19393 Segment
X19393 N19393 N19394 Segment
X19394 N19394 N19395 Segment
X19395 N19395 N19396 Segment
X19396 N19396 N19397 Segment
X19397 N19397 N19398 Segment
X19398 N19398 N19399 Segment
X19399 N19399 N19400 Segment
X19400 N19400 N19401 Segment
X19401 N19401 N19402 Segment
X19402 N19402 N19403 Segment
X19403 N19403 N19404 Segment
X19404 N19404 N19405 Segment
X19405 N19405 N19406 Segment
X19406 N19406 N19407 Segment
X19407 N19407 N19408 Segment
X19408 N19408 N19409 Segment
X19409 N19409 N19410 Segment
X19410 N19410 N19411 Segment
X19411 N19411 N19412 Segment
X19412 N19412 N19413 Segment
X19413 N19413 N19414 Segment
X19414 N19414 N19415 Segment
X19415 N19415 N19416 Segment
X19416 N19416 N19417 Segment
X19417 N19417 N19418 Segment
X19418 N19418 N19419 Segment
X19419 N19419 N19420 Segment
X19420 N19420 N19421 Segment
X19421 N19421 N19422 Segment
X19422 N19422 N19423 Segment
X19423 N19423 N19424 Segment
X19424 N19424 N19425 Segment
X19425 N19425 N19426 Segment
X19426 N19426 N19427 Segment
X19427 N19427 N19428 Segment
X19428 N19428 N19429 Segment
X19429 N19429 N19430 Segment
X19430 N19430 N19431 Segment
X19431 N19431 N19432 Segment
X19432 N19432 N19433 Segment
X19433 N19433 N19434 Segment
X19434 N19434 N19435 Segment
X19435 N19435 N19436 Segment
X19436 N19436 N19437 Segment
X19437 N19437 N19438 Segment
X19438 N19438 N19439 Segment
X19439 N19439 N19440 Segment
X19440 N19440 N19441 Segment
X19441 N19441 N19442 Segment
X19442 N19442 N19443 Segment
X19443 N19443 N19444 Segment
X19444 N19444 N19445 Segment
X19445 N19445 N19446 Segment
X19446 N19446 N19447 Segment
X19447 N19447 N19448 Segment
X19448 N19448 N19449 Segment
X19449 N19449 N19450 Segment
X19450 N19450 N19451 Segment
X19451 N19451 N19452 Segment
X19452 N19452 N19453 Segment
X19453 N19453 N19454 Segment
X19454 N19454 N19455 Segment
X19455 N19455 N19456 Segment
X19456 N19456 N19457 Segment
X19457 N19457 N19458 Segment
X19458 N19458 N19459 Segment
X19459 N19459 N19460 Segment
X19460 N19460 N19461 Segment
X19461 N19461 N19462 Segment
X19462 N19462 N19463 Segment
X19463 N19463 N19464 Segment
X19464 N19464 N19465 Segment
X19465 N19465 N19466 Segment
X19466 N19466 N19467 Segment
X19467 N19467 N19468 Segment
X19468 N19468 N19469 Segment
X19469 N19469 N19470 Segment
X19470 N19470 N19471 Segment
X19471 N19471 N19472 Segment
X19472 N19472 N19473 Segment
X19473 N19473 N19474 Segment
X19474 N19474 N19475 Segment
X19475 N19475 N19476 Segment
X19476 N19476 N19477 Segment
X19477 N19477 N19478 Segment
X19478 N19478 N19479 Segment
X19479 N19479 N19480 Segment
X19480 N19480 N19481 Segment
X19481 N19481 N19482 Segment
X19482 N19482 N19483 Segment
X19483 N19483 N19484 Segment
X19484 N19484 N19485 Segment
X19485 N19485 N19486 Segment
X19486 N19486 N19487 Segment
X19487 N19487 N19488 Segment
X19488 N19488 N19489 Segment
X19489 N19489 N19490 Segment
X19490 N19490 N19491 Segment
X19491 N19491 N19492 Segment
X19492 N19492 N19493 Segment
X19493 N19493 N19494 Segment
X19494 N19494 N19495 Segment
X19495 N19495 N19496 Segment
X19496 N19496 N19497 Segment
X19497 N19497 N19498 Segment
X19498 N19498 N19499 Segment
X19499 N19499 N19500 Segment
X19500 N19500 N19501 Segment
X19501 N19501 N19502 Segment
X19502 N19502 N19503 Segment
X19503 N19503 N19504 Segment
X19504 N19504 N19505 Segment
X19505 N19505 N19506 Segment
X19506 N19506 N19507 Segment
X19507 N19507 N19508 Segment
X19508 N19508 N19509 Segment
X19509 N19509 N19510 Segment
X19510 N19510 N19511 Segment
X19511 N19511 N19512 Segment
X19512 N19512 N19513 Segment
X19513 N19513 N19514 Segment
X19514 N19514 N19515 Segment
X19515 N19515 N19516 Segment
X19516 N19516 N19517 Segment
X19517 N19517 N19518 Segment
X19518 N19518 N19519 Segment
X19519 N19519 N19520 Segment
X19520 N19520 N19521 Segment
X19521 N19521 N19522 Segment
X19522 N19522 N19523 Segment
X19523 N19523 N19524 Segment
X19524 N19524 N19525 Segment
X19525 N19525 N19526 Segment
X19526 N19526 N19527 Segment
X19527 N19527 N19528 Segment
X19528 N19528 N19529 Segment
X19529 N19529 N19530 Segment
X19530 N19530 N19531 Segment
X19531 N19531 N19532 Segment
X19532 N19532 N19533 Segment
X19533 N19533 N19534 Segment
X19534 N19534 N19535 Segment
X19535 N19535 N19536 Segment
X19536 N19536 N19537 Segment
X19537 N19537 N19538 Segment
X19538 N19538 N19539 Segment
X19539 N19539 N19540 Segment
X19540 N19540 N19541 Segment
X19541 N19541 N19542 Segment
X19542 N19542 N19543 Segment
X19543 N19543 N19544 Segment
X19544 N19544 N19545 Segment
X19545 N19545 N19546 Segment
X19546 N19546 N19547 Segment
X19547 N19547 N19548 Segment
X19548 N19548 N19549 Segment
X19549 N19549 N19550 Segment
X19550 N19550 N19551 Segment
X19551 N19551 N19552 Segment
X19552 N19552 N19553 Segment
X19553 N19553 N19554 Segment
X19554 N19554 N19555 Segment
X19555 N19555 N19556 Segment
X19556 N19556 N19557 Segment
X19557 N19557 N19558 Segment
X19558 N19558 N19559 Segment
X19559 N19559 N19560 Segment
X19560 N19560 N19561 Segment
X19561 N19561 N19562 Segment
X19562 N19562 N19563 Segment
X19563 N19563 N19564 Segment
X19564 N19564 N19565 Segment
X19565 N19565 N19566 Segment
X19566 N19566 N19567 Segment
X19567 N19567 N19568 Segment
X19568 N19568 N19569 Segment
X19569 N19569 N19570 Segment
X19570 N19570 N19571 Segment
X19571 N19571 N19572 Segment
X19572 N19572 N19573 Segment
X19573 N19573 N19574 Segment
X19574 N19574 N19575 Segment
X19575 N19575 N19576 Segment
X19576 N19576 N19577 Segment
X19577 N19577 N19578 Segment
X19578 N19578 N19579 Segment
X19579 N19579 N19580 Segment
X19580 N19580 N19581 Segment
X19581 N19581 N19582 Segment
X19582 N19582 N19583 Segment
X19583 N19583 N19584 Segment
X19584 N19584 N19585 Segment
X19585 N19585 N19586 Segment
X19586 N19586 N19587 Segment
X19587 N19587 N19588 Segment
X19588 N19588 N19589 Segment
X19589 N19589 N19590 Segment
X19590 N19590 N19591 Segment
X19591 N19591 N19592 Segment
X19592 N19592 N19593 Segment
X19593 N19593 N19594 Segment
X19594 N19594 N19595 Segment
X19595 N19595 N19596 Segment
X19596 N19596 N19597 Segment
X19597 N19597 N19598 Segment
X19598 N19598 N19599 Segment
X19599 N19599 N19600 Segment
X19600 N19600 N19601 Segment
X19601 N19601 N19602 Segment
X19602 N19602 N19603 Segment
X19603 N19603 N19604 Segment
X19604 N19604 N19605 Segment
X19605 N19605 N19606 Segment
X19606 N19606 N19607 Segment
X19607 N19607 N19608 Segment
X19608 N19608 N19609 Segment
X19609 N19609 N19610 Segment
X19610 N19610 N19611 Segment
X19611 N19611 N19612 Segment
X19612 N19612 N19613 Segment
X19613 N19613 N19614 Segment
X19614 N19614 N19615 Segment
X19615 N19615 N19616 Segment
X19616 N19616 N19617 Segment
X19617 N19617 N19618 Segment
X19618 N19618 N19619 Segment
X19619 N19619 N19620 Segment
X19620 N19620 N19621 Segment
X19621 N19621 N19622 Segment
X19622 N19622 N19623 Segment
X19623 N19623 N19624 Segment
X19624 N19624 N19625 Segment
X19625 N19625 N19626 Segment
X19626 N19626 N19627 Segment
X19627 N19627 N19628 Segment
X19628 N19628 N19629 Segment
X19629 N19629 N19630 Segment
X19630 N19630 N19631 Segment
X19631 N19631 N19632 Segment
X19632 N19632 N19633 Segment
X19633 N19633 N19634 Segment
X19634 N19634 N19635 Segment
X19635 N19635 N19636 Segment
X19636 N19636 N19637 Segment
X19637 N19637 N19638 Segment
X19638 N19638 N19639 Segment
X19639 N19639 N19640 Segment
X19640 N19640 N19641 Segment
X19641 N19641 N19642 Segment
X19642 N19642 N19643 Segment
X19643 N19643 N19644 Segment
X19644 N19644 N19645 Segment
X19645 N19645 N19646 Segment
X19646 N19646 N19647 Segment
X19647 N19647 N19648 Segment
X19648 N19648 N19649 Segment
X19649 N19649 N19650 Segment
X19650 N19650 N19651 Segment
X19651 N19651 N19652 Segment
X19652 N19652 N19653 Segment
X19653 N19653 N19654 Segment
X19654 N19654 N19655 Segment
X19655 N19655 N19656 Segment
X19656 N19656 N19657 Segment
X19657 N19657 N19658 Segment
X19658 N19658 N19659 Segment
X19659 N19659 N19660 Segment
X19660 N19660 N19661 Segment
X19661 N19661 N19662 Segment
X19662 N19662 N19663 Segment
X19663 N19663 N19664 Segment
X19664 N19664 N19665 Segment
X19665 N19665 N19666 Segment
X19666 N19666 N19667 Segment
X19667 N19667 N19668 Segment
X19668 N19668 N19669 Segment
X19669 N19669 N19670 Segment
X19670 N19670 N19671 Segment
X19671 N19671 N19672 Segment
X19672 N19672 N19673 Segment
X19673 N19673 N19674 Segment
X19674 N19674 N19675 Segment
X19675 N19675 N19676 Segment
X19676 N19676 N19677 Segment
X19677 N19677 N19678 Segment
X19678 N19678 N19679 Segment
X19679 N19679 N19680 Segment
X19680 N19680 N19681 Segment
X19681 N19681 N19682 Segment
X19682 N19682 N19683 Segment
X19683 N19683 N19684 Segment
X19684 N19684 N19685 Segment
X19685 N19685 N19686 Segment
X19686 N19686 N19687 Segment
X19687 N19687 N19688 Segment
X19688 N19688 N19689 Segment
X19689 N19689 N19690 Segment
X19690 N19690 N19691 Segment
X19691 N19691 N19692 Segment
X19692 N19692 N19693 Segment
X19693 N19693 N19694 Segment
X19694 N19694 N19695 Segment
X19695 N19695 N19696 Segment
X19696 N19696 N19697 Segment
X19697 N19697 N19698 Segment
X19698 N19698 N19699 Segment
X19699 N19699 N19700 Segment
X19700 N19700 N19701 Segment
X19701 N19701 N19702 Segment
X19702 N19702 N19703 Segment
X19703 N19703 N19704 Segment
X19704 N19704 N19705 Segment
X19705 N19705 N19706 Segment
X19706 N19706 N19707 Segment
X19707 N19707 N19708 Segment
X19708 N19708 N19709 Segment
X19709 N19709 N19710 Segment
X19710 N19710 N19711 Segment
X19711 N19711 N19712 Segment
X19712 N19712 N19713 Segment
X19713 N19713 N19714 Segment
X19714 N19714 N19715 Segment
X19715 N19715 N19716 Segment
X19716 N19716 N19717 Segment
X19717 N19717 N19718 Segment
X19718 N19718 N19719 Segment
X19719 N19719 N19720 Segment
X19720 N19720 N19721 Segment
X19721 N19721 N19722 Segment
X19722 N19722 N19723 Segment
X19723 N19723 N19724 Segment
X19724 N19724 N19725 Segment
X19725 N19725 N19726 Segment
X19726 N19726 N19727 Segment
X19727 N19727 N19728 Segment
X19728 N19728 N19729 Segment
X19729 N19729 N19730 Segment
X19730 N19730 N19731 Segment
X19731 N19731 N19732 Segment
X19732 N19732 N19733 Segment
X19733 N19733 N19734 Segment
X19734 N19734 N19735 Segment
X19735 N19735 N19736 Segment
X19736 N19736 N19737 Segment
X19737 N19737 N19738 Segment
X19738 N19738 N19739 Segment
X19739 N19739 N19740 Segment
X19740 N19740 N19741 Segment
X19741 N19741 N19742 Segment
X19742 N19742 N19743 Segment
X19743 N19743 N19744 Segment
X19744 N19744 N19745 Segment
X19745 N19745 N19746 Segment
X19746 N19746 N19747 Segment
X19747 N19747 N19748 Segment
X19748 N19748 N19749 Segment
X19749 N19749 N19750 Segment
X19750 N19750 N19751 Segment
X19751 N19751 N19752 Segment
X19752 N19752 N19753 Segment
X19753 N19753 N19754 Segment
X19754 N19754 N19755 Segment
X19755 N19755 N19756 Segment
X19756 N19756 N19757 Segment
X19757 N19757 N19758 Segment
X19758 N19758 N19759 Segment
X19759 N19759 N19760 Segment
X19760 N19760 N19761 Segment
X19761 N19761 N19762 Segment
X19762 N19762 N19763 Segment
X19763 N19763 N19764 Segment
X19764 N19764 N19765 Segment
X19765 N19765 N19766 Segment
X19766 N19766 N19767 Segment
X19767 N19767 N19768 Segment
X19768 N19768 N19769 Segment
X19769 N19769 N19770 Segment
X19770 N19770 N19771 Segment
X19771 N19771 N19772 Segment
X19772 N19772 N19773 Segment
X19773 N19773 N19774 Segment
X19774 N19774 N19775 Segment
X19775 N19775 N19776 Segment
X19776 N19776 N19777 Segment
X19777 N19777 N19778 Segment
X19778 N19778 N19779 Segment
X19779 N19779 N19780 Segment
X19780 N19780 N19781 Segment
X19781 N19781 N19782 Segment
X19782 N19782 N19783 Segment
X19783 N19783 N19784 Segment
X19784 N19784 N19785 Segment
X19785 N19785 N19786 Segment
X19786 N19786 N19787 Segment
X19787 N19787 N19788 Segment
X19788 N19788 N19789 Segment
X19789 N19789 N19790 Segment
X19790 N19790 N19791 Segment
X19791 N19791 N19792 Segment
X19792 N19792 N19793 Segment
X19793 N19793 N19794 Segment
X19794 N19794 N19795 Segment
X19795 N19795 N19796 Segment
X19796 N19796 N19797 Segment
X19797 N19797 N19798 Segment
X19798 N19798 N19799 Segment
X19799 N19799 N19800 Segment
X19800 N19800 N19801 Segment
X19801 N19801 N19802 Segment
X19802 N19802 N19803 Segment
X19803 N19803 N19804 Segment
X19804 N19804 N19805 Segment
X19805 N19805 N19806 Segment
X19806 N19806 N19807 Segment
X19807 N19807 N19808 Segment
X19808 N19808 N19809 Segment
X19809 N19809 N19810 Segment
X19810 N19810 N19811 Segment
X19811 N19811 N19812 Segment
X19812 N19812 N19813 Segment
X19813 N19813 N19814 Segment
X19814 N19814 N19815 Segment
X19815 N19815 N19816 Segment
X19816 N19816 N19817 Segment
X19817 N19817 N19818 Segment
X19818 N19818 N19819 Segment
X19819 N19819 N19820 Segment
X19820 N19820 N19821 Segment
X19821 N19821 N19822 Segment
X19822 N19822 N19823 Segment
X19823 N19823 N19824 Segment
X19824 N19824 N19825 Segment
X19825 N19825 N19826 Segment
X19826 N19826 N19827 Segment
X19827 N19827 N19828 Segment
X19828 N19828 N19829 Segment
X19829 N19829 N19830 Segment
X19830 N19830 N19831 Segment
X19831 N19831 N19832 Segment
X19832 N19832 N19833 Segment
X19833 N19833 N19834 Segment
X19834 N19834 N19835 Segment
X19835 N19835 N19836 Segment
X19836 N19836 N19837 Segment
X19837 N19837 N19838 Segment
X19838 N19838 N19839 Segment
X19839 N19839 N19840 Segment
X19840 N19840 N19841 Segment
X19841 N19841 N19842 Segment
X19842 N19842 N19843 Segment
X19843 N19843 N19844 Segment
X19844 N19844 N19845 Segment
X19845 N19845 N19846 Segment
X19846 N19846 N19847 Segment
X19847 N19847 N19848 Segment
X19848 N19848 N19849 Segment
X19849 N19849 N19850 Segment
X19850 N19850 N19851 Segment
X19851 N19851 N19852 Segment
X19852 N19852 N19853 Segment
X19853 N19853 N19854 Segment
X19854 N19854 N19855 Segment
X19855 N19855 N19856 Segment
X19856 N19856 N19857 Segment
X19857 N19857 N19858 Segment
X19858 N19858 N19859 Segment
X19859 N19859 N19860 Segment
X19860 N19860 N19861 Segment
X19861 N19861 N19862 Segment
X19862 N19862 N19863 Segment
X19863 N19863 N19864 Segment
X19864 N19864 N19865 Segment
X19865 N19865 N19866 Segment
X19866 N19866 N19867 Segment
X19867 N19867 N19868 Segment
X19868 N19868 N19869 Segment
X19869 N19869 N19870 Segment
X19870 N19870 N19871 Segment
X19871 N19871 N19872 Segment
X19872 N19872 N19873 Segment
X19873 N19873 N19874 Segment
X19874 N19874 N19875 Segment
X19875 N19875 N19876 Segment
X19876 N19876 N19877 Segment
X19877 N19877 N19878 Segment
X19878 N19878 N19879 Segment
X19879 N19879 N19880 Segment
X19880 N19880 N19881 Segment
X19881 N19881 N19882 Segment
X19882 N19882 N19883 Segment
X19883 N19883 N19884 Segment
X19884 N19884 N19885 Segment
X19885 N19885 N19886 Segment
X19886 N19886 N19887 Segment
X19887 N19887 N19888 Segment
X19888 N19888 N19889 Segment
X19889 N19889 N19890 Segment
X19890 N19890 N19891 Segment
X19891 N19891 N19892 Segment
X19892 N19892 N19893 Segment
X19893 N19893 N19894 Segment
X19894 N19894 N19895 Segment
X19895 N19895 N19896 Segment
X19896 N19896 N19897 Segment
X19897 N19897 N19898 Segment
X19898 N19898 N19899 Segment
X19899 N19899 N19900 Segment
X19900 N19900 N19901 Segment
X19901 N19901 N19902 Segment
X19902 N19902 N19903 Segment
X19903 N19903 N19904 Segment
X19904 N19904 N19905 Segment
X19905 N19905 N19906 Segment
X19906 N19906 N19907 Segment
X19907 N19907 N19908 Segment
X19908 N19908 N19909 Segment
X19909 N19909 N19910 Segment
X19910 N19910 N19911 Segment
X19911 N19911 N19912 Segment
X19912 N19912 N19913 Segment
X19913 N19913 N19914 Segment
X19914 N19914 N19915 Segment
X19915 N19915 N19916 Segment
X19916 N19916 N19917 Segment
X19917 N19917 N19918 Segment
X19918 N19918 N19919 Segment
X19919 N19919 N19920 Segment
X19920 N19920 N19921 Segment
X19921 N19921 N19922 Segment
X19922 N19922 N19923 Segment
X19923 N19923 N19924 Segment
X19924 N19924 N19925 Segment
X19925 N19925 N19926 Segment
X19926 N19926 N19927 Segment
X19927 N19927 N19928 Segment
X19928 N19928 N19929 Segment
X19929 N19929 N19930 Segment
X19930 N19930 N19931 Segment
X19931 N19931 N19932 Segment
X19932 N19932 N19933 Segment
X19933 N19933 N19934 Segment
X19934 N19934 N19935 Segment
X19935 N19935 N19936 Segment
X19936 N19936 N19937 Segment
X19937 N19937 N19938 Segment
X19938 N19938 N19939 Segment
X19939 N19939 N19940 Segment
X19940 N19940 N19941 Segment
X19941 N19941 N19942 Segment
X19942 N19942 N19943 Segment
X19943 N19943 N19944 Segment
X19944 N19944 N19945 Segment
X19945 N19945 N19946 Segment
X19946 N19946 N19947 Segment
X19947 N19947 N19948 Segment
X19948 N19948 N19949 Segment
X19949 N19949 N19950 Segment
X19950 N19950 N19951 Segment
X19951 N19951 N19952 Segment
X19952 N19952 N19953 Segment
X19953 N19953 N19954 Segment
X19954 N19954 N19955 Segment
X19955 N19955 N19956 Segment
X19956 N19956 N19957 Segment
X19957 N19957 N19958 Segment
X19958 N19958 N19959 Segment
X19959 N19959 N19960 Segment
X19960 N19960 N19961 Segment
X19961 N19961 N19962 Segment
X19962 N19962 N19963 Segment
X19963 N19963 N19964 Segment
X19964 N19964 N19965 Segment
X19965 N19965 N19966 Segment
X19966 N19966 N19967 Segment
X19967 N19967 N19968 Segment
X19968 N19968 N19969 Segment
X19969 N19969 N19970 Segment
X19970 N19970 N19971 Segment
X19971 N19971 N19972 Segment
X19972 N19972 N19973 Segment
X19973 N19973 N19974 Segment
X19974 N19974 N19975 Segment
X19975 N19975 N19976 Segment
X19976 N19976 N19977 Segment
X19977 N19977 N19978 Segment
X19978 N19978 N19979 Segment
X19979 N19979 N19980 Segment
X19980 N19980 N19981 Segment
X19981 N19981 N19982 Segment
X19982 N19982 N19983 Segment
X19983 N19983 N19984 Segment
X19984 N19984 N19985 Segment
X19985 N19985 N19986 Segment
X19986 N19986 N19987 Segment
X19987 N19987 N19988 Segment
X19988 N19988 N19989 Segment
X19989 N19989 N19990 Segment
X19990 N19990 N19991 Segment
X19991 N19991 N19992 Segment
X19992 N19992 N19993 Segment
X19993 N19993 N19994 Segment
X19994 N19994 N19995 Segment
X19995 N19995 N19996 Segment
X19996 N19996 N19997 Segment
X19997 N19997 N19998 Segment
X19998 N19998 N19999 Segment
X19999 N19999 N20000 Segment
X20000 N20000 N20001 Segment
X20001 N20001 N20002 Segment
X20002 N20002 N20003 Segment
X20003 N20003 N20004 Segment
X20004 N20004 N20005 Segment
X20005 N20005 N20006 Segment
X20006 N20006 N20007 Segment
X20007 N20007 N20008 Segment
X20008 N20008 N20009 Segment
X20009 N20009 N20010 Segment
X20010 N20010 N20011 Segment
X20011 N20011 N20012 Segment
X20012 N20012 N20013 Segment
X20013 N20013 N20014 Segment
X20014 N20014 N20015 Segment
X20015 N20015 N20016 Segment
X20016 N20016 N20017 Segment
X20017 N20017 N20018 Segment
X20018 N20018 N20019 Segment
X20019 N20019 N20020 Segment
X20020 N20020 N20021 Segment
X20021 N20021 N20022 Segment
X20022 N20022 N20023 Segment
X20023 N20023 N20024 Segment
X20024 N20024 N20025 Segment
X20025 N20025 N20026 Segment
X20026 N20026 N20027 Segment
X20027 N20027 N20028 Segment
X20028 N20028 N20029 Segment
X20029 N20029 N20030 Segment
X20030 N20030 N20031 Segment
X20031 N20031 N20032 Segment
X20032 N20032 N20033 Segment
X20033 N20033 N20034 Segment
X20034 N20034 N20035 Segment
X20035 N20035 N20036 Segment
X20036 N20036 N20037 Segment
X20037 N20037 N20038 Segment
X20038 N20038 N20039 Segment
X20039 N20039 N20040 Segment
X20040 N20040 N20041 Segment
X20041 N20041 N20042 Segment
X20042 N20042 N20043 Segment
X20043 N20043 N20044 Segment
X20044 N20044 N20045 Segment
X20045 N20045 N20046 Segment
X20046 N20046 N20047 Segment
X20047 N20047 N20048 Segment
X20048 N20048 N20049 Segment
X20049 N20049 N20050 Segment
X20050 N20050 N20051 Segment
X20051 N20051 N20052 Segment
X20052 N20052 N20053 Segment
X20053 N20053 N20054 Segment
X20054 N20054 N20055 Segment
X20055 N20055 N20056 Segment
X20056 N20056 N20057 Segment
X20057 N20057 N20058 Segment
X20058 N20058 N20059 Segment
X20059 N20059 N20060 Segment
X20060 N20060 N20061 Segment
X20061 N20061 N20062 Segment
X20062 N20062 N20063 Segment
X20063 N20063 N20064 Segment
X20064 N20064 N20065 Segment
X20065 N20065 N20066 Segment
X20066 N20066 N20067 Segment
X20067 N20067 N20068 Segment
X20068 N20068 N20069 Segment
X20069 N20069 N20070 Segment
X20070 N20070 N20071 Segment
X20071 N20071 N20072 Segment
X20072 N20072 N20073 Segment
X20073 N20073 N20074 Segment
X20074 N20074 N20075 Segment
X20075 N20075 N20076 Segment
X20076 N20076 N20077 Segment
X20077 N20077 N20078 Segment
X20078 N20078 N20079 Segment
X20079 N20079 N20080 Segment
X20080 N20080 N20081 Segment
X20081 N20081 N20082 Segment
X20082 N20082 N20083 Segment
X20083 N20083 N20084 Segment
X20084 N20084 N20085 Segment
X20085 N20085 N20086 Segment
X20086 N20086 N20087 Segment
X20087 N20087 N20088 Segment
X20088 N20088 N20089 Segment
X20089 N20089 N20090 Segment
X20090 N20090 N20091 Segment
X20091 N20091 N20092 Segment
X20092 N20092 N20093 Segment
X20093 N20093 N20094 Segment
X20094 N20094 N20095 Segment
X20095 N20095 N20096 Segment
X20096 N20096 N20097 Segment
X20097 N20097 N20098 Segment
X20098 N20098 N20099 Segment
X20099 N20099 N20100 Segment
X20100 N20100 N20101 Segment
X20101 N20101 N20102 Segment
X20102 N20102 N20103 Segment
X20103 N20103 N20104 Segment
X20104 N20104 N20105 Segment
X20105 N20105 N20106 Segment
X20106 N20106 N20107 Segment
X20107 N20107 N20108 Segment
X20108 N20108 N20109 Segment
X20109 N20109 N20110 Segment
X20110 N20110 N20111 Segment
X20111 N20111 N20112 Segment
X20112 N20112 N20113 Segment
X20113 N20113 N20114 Segment
X20114 N20114 N20115 Segment
X20115 N20115 N20116 Segment
X20116 N20116 N20117 Segment
X20117 N20117 N20118 Segment
X20118 N20118 N20119 Segment
X20119 N20119 N20120 Segment
X20120 N20120 N20121 Segment
X20121 N20121 N20122 Segment
X20122 N20122 N20123 Segment
X20123 N20123 N20124 Segment
X20124 N20124 N20125 Segment
X20125 N20125 N20126 Segment
X20126 N20126 N20127 Segment
X20127 N20127 N20128 Segment
X20128 N20128 N20129 Segment
X20129 N20129 N20130 Segment
X20130 N20130 N20131 Segment
X20131 N20131 N20132 Segment
X20132 N20132 N20133 Segment
X20133 N20133 N20134 Segment
X20134 N20134 N20135 Segment
X20135 N20135 N20136 Segment
X20136 N20136 N20137 Segment
X20137 N20137 N20138 Segment
X20138 N20138 N20139 Segment
X20139 N20139 N20140 Segment
X20140 N20140 N20141 Segment
X20141 N20141 N20142 Segment
X20142 N20142 N20143 Segment
X20143 N20143 N20144 Segment
X20144 N20144 N20145 Segment
X20145 N20145 N20146 Segment
X20146 N20146 N20147 Segment
X20147 N20147 N20148 Segment
X20148 N20148 N20149 Segment
X20149 N20149 N20150 Segment
X20150 N20150 N20151 Segment
X20151 N20151 N20152 Segment
X20152 N20152 N20153 Segment
X20153 N20153 N20154 Segment
X20154 N20154 N20155 Segment
X20155 N20155 N20156 Segment
X20156 N20156 N20157 Segment
X20157 N20157 N20158 Segment
X20158 N20158 N20159 Segment
X20159 N20159 N20160 Segment
X20160 N20160 N20161 Segment
X20161 N20161 N20162 Segment
X20162 N20162 N20163 Segment
X20163 N20163 N20164 Segment
X20164 N20164 N20165 Segment
X20165 N20165 N20166 Segment
X20166 N20166 N20167 Segment
X20167 N20167 N20168 Segment
X20168 N20168 N20169 Segment
X20169 N20169 N20170 Segment
X20170 N20170 N20171 Segment
X20171 N20171 N20172 Segment
X20172 N20172 N20173 Segment
X20173 N20173 N20174 Segment
X20174 N20174 N20175 Segment
X20175 N20175 N20176 Segment
X20176 N20176 N20177 Segment
X20177 N20177 N20178 Segment
X20178 N20178 N20179 Segment
X20179 N20179 N20180 Segment
X20180 N20180 N20181 Segment
X20181 N20181 N20182 Segment
X20182 N20182 N20183 Segment
X20183 N20183 N20184 Segment
X20184 N20184 N20185 Segment
X20185 N20185 N20186 Segment
X20186 N20186 N20187 Segment
X20187 N20187 N20188 Segment
X20188 N20188 N20189 Segment
X20189 N20189 N20190 Segment
X20190 N20190 N20191 Segment
X20191 N20191 N20192 Segment
X20192 N20192 N20193 Segment
X20193 N20193 N20194 Segment
X20194 N20194 N20195 Segment
X20195 N20195 N20196 Segment
X20196 N20196 N20197 Segment
X20197 N20197 N20198 Segment
X20198 N20198 N20199 Segment
X20199 N20199 N20200 Segment
X20200 N20200 N20201 Segment
X20201 N20201 N20202 Segment
X20202 N20202 N20203 Segment
X20203 N20203 N20204 Segment
X20204 N20204 N20205 Segment
X20205 N20205 N20206 Segment
X20206 N20206 N20207 Segment
X20207 N20207 N20208 Segment
X20208 N20208 N20209 Segment
X20209 N20209 N20210 Segment
X20210 N20210 N20211 Segment
X20211 N20211 N20212 Segment
X20212 N20212 N20213 Segment
X20213 N20213 N20214 Segment
X20214 N20214 N20215 Segment
X20215 N20215 N20216 Segment
X20216 N20216 N20217 Segment
X20217 N20217 N20218 Segment
X20218 N20218 N20219 Segment
X20219 N20219 N20220 Segment
X20220 N20220 N20221 Segment
X20221 N20221 N20222 Segment
X20222 N20222 N20223 Segment
X20223 N20223 N20224 Segment
X20224 N20224 N20225 Segment
X20225 N20225 N20226 Segment
X20226 N20226 N20227 Segment
X20227 N20227 N20228 Segment
X20228 N20228 N20229 Segment
X20229 N20229 N20230 Segment
X20230 N20230 N20231 Segment
X20231 N20231 N20232 Segment
X20232 N20232 N20233 Segment
X20233 N20233 N20234 Segment
X20234 N20234 N20235 Segment
X20235 N20235 N20236 Segment
X20236 N20236 N20237 Segment
X20237 N20237 N20238 Segment
X20238 N20238 N20239 Segment
X20239 N20239 N20240 Segment
X20240 N20240 N20241 Segment
X20241 N20241 N20242 Segment
X20242 N20242 N20243 Segment
X20243 N20243 N20244 Segment
X20244 N20244 N20245 Segment
X20245 N20245 N20246 Segment
X20246 N20246 N20247 Segment
X20247 N20247 N20248 Segment
X20248 N20248 N20249 Segment
X20249 N20249 N20250 Segment
X20250 N20250 N20251 Segment
X20251 N20251 N20252 Segment
X20252 N20252 N20253 Segment
X20253 N20253 N20254 Segment
X20254 N20254 N20255 Segment
X20255 N20255 N20256 Segment
X20256 N20256 N20257 Segment
X20257 N20257 N20258 Segment
X20258 N20258 N20259 Segment
X20259 N20259 N20260 Segment
X20260 N20260 N20261 Segment
X20261 N20261 N20262 Segment
X20262 N20262 N20263 Segment
X20263 N20263 N20264 Segment
X20264 N20264 N20265 Segment
X20265 N20265 N20266 Segment
X20266 N20266 N20267 Segment
X20267 N20267 N20268 Segment
X20268 N20268 N20269 Segment
X20269 N20269 N20270 Segment
X20270 N20270 N20271 Segment
X20271 N20271 N20272 Segment
X20272 N20272 N20273 Segment
X20273 N20273 N20274 Segment
X20274 N20274 N20275 Segment
X20275 N20275 N20276 Segment
X20276 N20276 N20277 Segment
X20277 N20277 N20278 Segment
X20278 N20278 N20279 Segment
X20279 N20279 N20280 Segment
X20280 N20280 N20281 Segment
X20281 N20281 N20282 Segment
X20282 N20282 N20283 Segment
X20283 N20283 N20284 Segment
X20284 N20284 N20285 Segment
X20285 N20285 N20286 Segment
X20286 N20286 N20287 Segment
X20287 N20287 N20288 Segment
X20288 N20288 N20289 Segment
X20289 N20289 N20290 Segment
X20290 N20290 N20291 Segment
X20291 N20291 N20292 Segment
X20292 N20292 N20293 Segment
X20293 N20293 N20294 Segment
X20294 N20294 N20295 Segment
X20295 N20295 N20296 Segment
X20296 N20296 N20297 Segment
X20297 N20297 N20298 Segment
X20298 N20298 N20299 Segment
X20299 N20299 N20300 Segment
X20300 N20300 N20301 Segment
X20301 N20301 N20302 Segment
X20302 N20302 N20303 Segment
X20303 N20303 N20304 Segment
X20304 N20304 N20305 Segment
X20305 N20305 N20306 Segment
X20306 N20306 N20307 Segment
X20307 N20307 N20308 Segment
X20308 N20308 N20309 Segment
X20309 N20309 N20310 Segment
X20310 N20310 N20311 Segment
X20311 N20311 N20312 Segment
X20312 N20312 N20313 Segment
X20313 N20313 N20314 Segment
X20314 N20314 N20315 Segment
X20315 N20315 N20316 Segment
X20316 N20316 N20317 Segment
X20317 N20317 N20318 Segment
X20318 N20318 N20319 Segment
X20319 N20319 N20320 Segment
X20320 N20320 N20321 Segment
X20321 N20321 N20322 Segment
X20322 N20322 N20323 Segment
X20323 N20323 N20324 Segment
X20324 N20324 N20325 Segment
X20325 N20325 N20326 Segment
X20326 N20326 N20327 Segment
X20327 N20327 N20328 Segment
X20328 N20328 N20329 Segment
X20329 N20329 N20330 Segment
X20330 N20330 N20331 Segment
X20331 N20331 N20332 Segment
X20332 N20332 N20333 Segment
X20333 N20333 N20334 Segment
X20334 N20334 N20335 Segment
X20335 N20335 N20336 Segment
X20336 N20336 N20337 Segment
X20337 N20337 N20338 Segment
X20338 N20338 N20339 Segment
X20339 N20339 N20340 Segment
X20340 N20340 N20341 Segment
X20341 N20341 N20342 Segment
X20342 N20342 N20343 Segment
X20343 N20343 N20344 Segment
X20344 N20344 N20345 Segment
X20345 N20345 N20346 Segment
X20346 N20346 N20347 Segment
X20347 N20347 N20348 Segment
X20348 N20348 N20349 Segment
X20349 N20349 N20350 Segment
X20350 N20350 N20351 Segment
X20351 N20351 N20352 Segment
X20352 N20352 N20353 Segment
X20353 N20353 N20354 Segment
X20354 N20354 N20355 Segment
X20355 N20355 N20356 Segment
X20356 N20356 N20357 Segment
X20357 N20357 N20358 Segment
X20358 N20358 N20359 Segment
X20359 N20359 N20360 Segment
X20360 N20360 N20361 Segment
X20361 N20361 N20362 Segment
X20362 N20362 N20363 Segment
X20363 N20363 N20364 Segment
X20364 N20364 N20365 Segment
X20365 N20365 N20366 Segment
X20366 N20366 N20367 Segment
X20367 N20367 N20368 Segment
X20368 N20368 N20369 Segment
X20369 N20369 N20370 Segment
X20370 N20370 N20371 Segment
X20371 N20371 N20372 Segment
X20372 N20372 N20373 Segment
X20373 N20373 N20374 Segment
X20374 N20374 N20375 Segment
X20375 N20375 N20376 Segment
X20376 N20376 N20377 Segment
X20377 N20377 N20378 Segment
X20378 N20378 N20379 Segment
X20379 N20379 N20380 Segment
X20380 N20380 N20381 Segment
X20381 N20381 N20382 Segment
X20382 N20382 N20383 Segment
X20383 N20383 N20384 Segment
X20384 N20384 N20385 Segment
X20385 N20385 N20386 Segment
X20386 N20386 N20387 Segment
X20387 N20387 N20388 Segment
X20388 N20388 N20389 Segment
X20389 N20389 N20390 Segment
X20390 N20390 N20391 Segment
X20391 N20391 N20392 Segment
X20392 N20392 N20393 Segment
X20393 N20393 N20394 Segment
X20394 N20394 N20395 Segment
X20395 N20395 N20396 Segment
X20396 N20396 N20397 Segment
X20397 N20397 N20398 Segment
X20398 N20398 N20399 Segment
X20399 N20399 N20400 Segment
X20400 N20400 N20401 Segment
X20401 N20401 N20402 Segment
X20402 N20402 N20403 Segment
X20403 N20403 N20404 Segment
X20404 N20404 N20405 Segment
X20405 N20405 N20406 Segment
X20406 N20406 N20407 Segment
X20407 N20407 N20408 Segment
X20408 N20408 N20409 Segment
X20409 N20409 N20410 Segment
X20410 N20410 N20411 Segment
X20411 N20411 N20412 Segment
X20412 N20412 N20413 Segment
X20413 N20413 N20414 Segment
X20414 N20414 N20415 Segment
X20415 N20415 N20416 Segment
X20416 N20416 N20417 Segment
X20417 N20417 N20418 Segment
X20418 N20418 N20419 Segment
X20419 N20419 N20420 Segment
X20420 N20420 N20421 Segment
X20421 N20421 N20422 Segment
X20422 N20422 N20423 Segment
X20423 N20423 N20424 Segment
X20424 N20424 N20425 Segment
X20425 N20425 N20426 Segment
X20426 N20426 N20427 Segment
X20427 N20427 N20428 Segment
X20428 N20428 N20429 Segment
X20429 N20429 N20430 Segment
X20430 N20430 N20431 Segment
X20431 N20431 N20432 Segment
X20432 N20432 N20433 Segment
X20433 N20433 N20434 Segment
X20434 N20434 N20435 Segment
X20435 N20435 N20436 Segment
X20436 N20436 N20437 Segment
X20437 N20437 N20438 Segment
X20438 N20438 N20439 Segment
X20439 N20439 N20440 Segment
X20440 N20440 N20441 Segment
X20441 N20441 N20442 Segment
X20442 N20442 N20443 Segment
X20443 N20443 N20444 Segment
X20444 N20444 N20445 Segment
X20445 N20445 N20446 Segment
X20446 N20446 N20447 Segment
X20447 N20447 N20448 Segment
X20448 N20448 N20449 Segment
X20449 N20449 N20450 Segment
X20450 N20450 N20451 Segment
X20451 N20451 N20452 Segment
X20452 N20452 N20453 Segment
X20453 N20453 N20454 Segment
X20454 N20454 N20455 Segment
X20455 N20455 N20456 Segment
X20456 N20456 N20457 Segment
X20457 N20457 N20458 Segment
X20458 N20458 N20459 Segment
X20459 N20459 N20460 Segment
X20460 N20460 N20461 Segment
X20461 N20461 N20462 Segment
X20462 N20462 N20463 Segment
X20463 N20463 N20464 Segment
X20464 N20464 N20465 Segment
X20465 N20465 N20466 Segment
X20466 N20466 N20467 Segment
X20467 N20467 N20468 Segment
X20468 N20468 N20469 Segment
X20469 N20469 N20470 Segment
X20470 N20470 N20471 Segment
X20471 N20471 N20472 Segment
X20472 N20472 N20473 Segment
X20473 N20473 N20474 Segment
X20474 N20474 N20475 Segment
X20475 N20475 N20476 Segment
X20476 N20476 N20477 Segment
X20477 N20477 N20478 Segment
X20478 N20478 N20479 Segment
X20479 N20479 N20480 Segment
X20480 N20480 N20481 Segment
X20481 N20481 N20482 Segment
X20482 N20482 N20483 Segment
X20483 N20483 N20484 Segment
X20484 N20484 N20485 Segment
X20485 N20485 N20486 Segment
X20486 N20486 N20487 Segment
X20487 N20487 N20488 Segment
X20488 N20488 N20489 Segment
X20489 N20489 N20490 Segment
X20490 N20490 N20491 Segment
X20491 N20491 N20492 Segment
X20492 N20492 N20493 Segment
X20493 N20493 N20494 Segment
X20494 N20494 N20495 Segment
X20495 N20495 N20496 Segment
X20496 N20496 N20497 Segment
X20497 N20497 N20498 Segment
X20498 N20498 N20499 Segment
X20499 N20499 N20500 Segment
X20500 N20500 N20501 Segment
X20501 N20501 N20502 Segment
X20502 N20502 N20503 Segment
X20503 N20503 N20504 Segment
X20504 N20504 N20505 Segment
X20505 N20505 N20506 Segment
X20506 N20506 N20507 Segment
X20507 N20507 N20508 Segment
X20508 N20508 N20509 Segment
X20509 N20509 N20510 Segment
X20510 N20510 N20511 Segment
X20511 N20511 N20512 Segment
X20512 N20512 N20513 Segment
X20513 N20513 N20514 Segment
X20514 N20514 N20515 Segment
X20515 N20515 N20516 Segment
X20516 N20516 N20517 Segment
X20517 N20517 N20518 Segment
X20518 N20518 N20519 Segment
X20519 N20519 N20520 Segment
X20520 N20520 N20521 Segment
X20521 N20521 N20522 Segment
X20522 N20522 N20523 Segment
X20523 N20523 N20524 Segment
X20524 N20524 N20525 Segment
X20525 N20525 N20526 Segment
X20526 N20526 N20527 Segment
X20527 N20527 N20528 Segment
X20528 N20528 N20529 Segment
X20529 N20529 N20530 Segment
X20530 N20530 N20531 Segment
X20531 N20531 N20532 Segment
X20532 N20532 N20533 Segment
X20533 N20533 N20534 Segment
X20534 N20534 N20535 Segment
X20535 N20535 N20536 Segment
X20536 N20536 N20537 Segment
X20537 N20537 N20538 Segment
X20538 N20538 N20539 Segment
X20539 N20539 N20540 Segment
X20540 N20540 N20541 Segment
X20541 N20541 N20542 Segment
X20542 N20542 N20543 Segment
X20543 N20543 N20544 Segment
X20544 N20544 N20545 Segment
X20545 N20545 N20546 Segment
X20546 N20546 N20547 Segment
X20547 N20547 N20548 Segment
X20548 N20548 N20549 Segment
X20549 N20549 N20550 Segment
X20550 N20550 N20551 Segment
X20551 N20551 N20552 Segment
X20552 N20552 N20553 Segment
X20553 N20553 N20554 Segment
X20554 N20554 N20555 Segment
X20555 N20555 N20556 Segment
X20556 N20556 N20557 Segment
X20557 N20557 N20558 Segment
X20558 N20558 N20559 Segment
X20559 N20559 N20560 Segment
X20560 N20560 N20561 Segment
X20561 N20561 N20562 Segment
X20562 N20562 N20563 Segment
X20563 N20563 N20564 Segment
X20564 N20564 N20565 Segment
X20565 N20565 N20566 Segment
X20566 N20566 N20567 Segment
X20567 N20567 N20568 Segment
X20568 N20568 N20569 Segment
X20569 N20569 N20570 Segment
X20570 N20570 N20571 Segment
X20571 N20571 N20572 Segment
X20572 N20572 N20573 Segment
X20573 N20573 N20574 Segment
X20574 N20574 N20575 Segment
X20575 N20575 N20576 Segment
X20576 N20576 N20577 Segment
X20577 N20577 N20578 Segment
X20578 N20578 N20579 Segment
X20579 N20579 N20580 Segment
X20580 N20580 N20581 Segment
X20581 N20581 N20582 Segment
X20582 N20582 N20583 Segment
X20583 N20583 N20584 Segment
X20584 N20584 N20585 Segment
X20585 N20585 N20586 Segment
X20586 N20586 N20587 Segment
X20587 N20587 N20588 Segment
X20588 N20588 N20589 Segment
X20589 N20589 N20590 Segment
X20590 N20590 N20591 Segment
X20591 N20591 N20592 Segment
X20592 N20592 N20593 Segment
X20593 N20593 N20594 Segment
X20594 N20594 N20595 Segment
X20595 N20595 N20596 Segment
X20596 N20596 N20597 Segment
X20597 N20597 N20598 Segment
X20598 N20598 N20599 Segment
X20599 N20599 N20600 Segment
X20600 N20600 N20601 Segment
X20601 N20601 N20602 Segment
X20602 N20602 N20603 Segment
X20603 N20603 N20604 Segment
X20604 N20604 N20605 Segment
X20605 N20605 N20606 Segment
X20606 N20606 N20607 Segment
X20607 N20607 N20608 Segment
X20608 N20608 N20609 Segment
X20609 N20609 N20610 Segment
X20610 N20610 N20611 Segment
X20611 N20611 N20612 Segment
X20612 N20612 N20613 Segment
X20613 N20613 N20614 Segment
X20614 N20614 N20615 Segment
X20615 N20615 N20616 Segment
X20616 N20616 N20617 Segment
X20617 N20617 N20618 Segment
X20618 N20618 N20619 Segment
X20619 N20619 N20620 Segment
X20620 N20620 N20621 Segment
X20621 N20621 N20622 Segment
X20622 N20622 N20623 Segment
X20623 N20623 N20624 Segment
X20624 N20624 N20625 Segment
X20625 N20625 N20626 Segment
X20626 N20626 N20627 Segment
X20627 N20627 N20628 Segment
X20628 N20628 N20629 Segment
X20629 N20629 N20630 Segment
X20630 N20630 N20631 Segment
X20631 N20631 N20632 Segment
X20632 N20632 N20633 Segment
X20633 N20633 N20634 Segment
X20634 N20634 N20635 Segment
X20635 N20635 N20636 Segment
X20636 N20636 N20637 Segment
X20637 N20637 N20638 Segment
X20638 N20638 N20639 Segment
X20639 N20639 N20640 Segment
X20640 N20640 N20641 Segment
X20641 N20641 N20642 Segment
X20642 N20642 N20643 Segment
X20643 N20643 N20644 Segment
X20644 N20644 N20645 Segment
X20645 N20645 N20646 Segment
X20646 N20646 N20647 Segment
X20647 N20647 N20648 Segment
X20648 N20648 N20649 Segment
X20649 N20649 N20650 Segment
X20650 N20650 N20651 Segment
X20651 N20651 N20652 Segment
X20652 N20652 N20653 Segment
X20653 N20653 N20654 Segment
X20654 N20654 N20655 Segment
X20655 N20655 N20656 Segment
X20656 N20656 N20657 Segment
X20657 N20657 N20658 Segment
X20658 N20658 N20659 Segment
X20659 N20659 N20660 Segment
X20660 N20660 N20661 Segment
X20661 N20661 N20662 Segment
X20662 N20662 N20663 Segment
X20663 N20663 N20664 Segment
X20664 N20664 N20665 Segment
X20665 N20665 N20666 Segment
X20666 N20666 N20667 Segment
X20667 N20667 N20668 Segment
X20668 N20668 N20669 Segment
X20669 N20669 N20670 Segment
X20670 N20670 N20671 Segment
X20671 N20671 N20672 Segment
X20672 N20672 N20673 Segment
X20673 N20673 N20674 Segment
X20674 N20674 N20675 Segment
X20675 N20675 N20676 Segment
X20676 N20676 N20677 Segment
X20677 N20677 N20678 Segment
X20678 N20678 N20679 Segment
X20679 N20679 N20680 Segment
X20680 N20680 N20681 Segment
X20681 N20681 N20682 Segment
X20682 N20682 N20683 Segment
X20683 N20683 N20684 Segment
X20684 N20684 N20685 Segment
X20685 N20685 N20686 Segment
X20686 N20686 N20687 Segment
X20687 N20687 N20688 Segment
X20688 N20688 N20689 Segment
X20689 N20689 N20690 Segment
X20690 N20690 N20691 Segment
X20691 N20691 N20692 Segment
X20692 N20692 N20693 Segment
X20693 N20693 N20694 Segment
X20694 N20694 N20695 Segment
X20695 N20695 N20696 Segment
X20696 N20696 N20697 Segment
X20697 N20697 N20698 Segment
X20698 N20698 N20699 Segment
X20699 N20699 N20700 Segment
X20700 N20700 N20701 Segment
X20701 N20701 N20702 Segment
X20702 N20702 N20703 Segment
X20703 N20703 N20704 Segment
X20704 N20704 N20705 Segment
X20705 N20705 N20706 Segment
X20706 N20706 N20707 Segment
X20707 N20707 N20708 Segment
X20708 N20708 N20709 Segment
X20709 N20709 N20710 Segment
X20710 N20710 N20711 Segment
X20711 N20711 N20712 Segment
X20712 N20712 N20713 Segment
X20713 N20713 N20714 Segment
X20714 N20714 N20715 Segment
X20715 N20715 N20716 Segment
X20716 N20716 N20717 Segment
X20717 N20717 N20718 Segment
X20718 N20718 N20719 Segment
X20719 N20719 N20720 Segment
X20720 N20720 N20721 Segment
X20721 N20721 N20722 Segment
X20722 N20722 N20723 Segment
X20723 N20723 N20724 Segment
X20724 N20724 N20725 Segment
X20725 N20725 N20726 Segment
X20726 N20726 N20727 Segment
X20727 N20727 N20728 Segment
X20728 N20728 N20729 Segment
X20729 N20729 N20730 Segment
X20730 N20730 N20731 Segment
X20731 N20731 N20732 Segment
X20732 N20732 N20733 Segment
X20733 N20733 N20734 Segment
X20734 N20734 N20735 Segment
X20735 N20735 N20736 Segment
X20736 N20736 N20737 Segment
X20737 N20737 N20738 Segment
X20738 N20738 N20739 Segment
X20739 N20739 N20740 Segment
X20740 N20740 N20741 Segment
X20741 N20741 N20742 Segment
X20742 N20742 N20743 Segment
X20743 N20743 N20744 Segment
X20744 N20744 N20745 Segment
X20745 N20745 N20746 Segment
X20746 N20746 N20747 Segment
X20747 N20747 N20748 Segment
X20748 N20748 N20749 Segment
X20749 N20749 N20750 Segment
X20750 N20750 N20751 Segment
X20751 N20751 N20752 Segment
X20752 N20752 N20753 Segment
X20753 N20753 N20754 Segment
X20754 N20754 N20755 Segment
X20755 N20755 N20756 Segment
X20756 N20756 N20757 Segment
X20757 N20757 N20758 Segment
X20758 N20758 N20759 Segment
X20759 N20759 N20760 Segment
X20760 N20760 N20761 Segment
X20761 N20761 N20762 Segment
X20762 N20762 N20763 Segment
X20763 N20763 N20764 Segment
X20764 N20764 N20765 Segment
X20765 N20765 N20766 Segment
X20766 N20766 N20767 Segment
X20767 N20767 N20768 Segment
X20768 N20768 N20769 Segment
X20769 N20769 N20770 Segment
X20770 N20770 N20771 Segment
X20771 N20771 N20772 Segment
X20772 N20772 N20773 Segment
X20773 N20773 N20774 Segment
X20774 N20774 N20775 Segment
X20775 N20775 N20776 Segment
X20776 N20776 N20777 Segment
X20777 N20777 N20778 Segment
X20778 N20778 N20779 Segment
X20779 N20779 N20780 Segment
X20780 N20780 N20781 Segment
X20781 N20781 N20782 Segment
X20782 N20782 N20783 Segment
X20783 N20783 N20784 Segment
X20784 N20784 N20785 Segment
X20785 N20785 N20786 Segment
X20786 N20786 N20787 Segment
X20787 N20787 N20788 Segment
X20788 N20788 N20789 Segment
X20789 N20789 N20790 Segment
X20790 N20790 N20791 Segment
X20791 N20791 N20792 Segment
X20792 N20792 N20793 Segment
X20793 N20793 N20794 Segment
X20794 N20794 N20795 Segment
X20795 N20795 N20796 Segment
X20796 N20796 N20797 Segment
X20797 N20797 N20798 Segment
X20798 N20798 N20799 Segment
X20799 N20799 N20800 Segment
X20800 N20800 N20801 Segment
X20801 N20801 N20802 Segment
X20802 N20802 N20803 Segment
X20803 N20803 N20804 Segment
X20804 N20804 N20805 Segment
X20805 N20805 N20806 Segment
X20806 N20806 N20807 Segment
X20807 N20807 N20808 Segment
X20808 N20808 N20809 Segment
X20809 N20809 N20810 Segment
X20810 N20810 N20811 Segment
X20811 N20811 N20812 Segment
X20812 N20812 N20813 Segment
X20813 N20813 N20814 Segment
X20814 N20814 N20815 Segment
X20815 N20815 N20816 Segment
X20816 N20816 N20817 Segment
X20817 N20817 N20818 Segment
X20818 N20818 N20819 Segment
X20819 N20819 N20820 Segment
X20820 N20820 N20821 Segment
X20821 N20821 N20822 Segment
X20822 N20822 N20823 Segment
X20823 N20823 N20824 Segment
X20824 N20824 N20825 Segment
X20825 N20825 N20826 Segment
X20826 N20826 N20827 Segment
X20827 N20827 N20828 Segment
X20828 N20828 N20829 Segment
X20829 N20829 N20830 Segment
X20830 N20830 N20831 Segment
X20831 N20831 N20832 Segment
X20832 N20832 N20833 Segment
X20833 N20833 N20834 Segment
X20834 N20834 N20835 Segment
X20835 N20835 N20836 Segment
X20836 N20836 N20837 Segment
X20837 N20837 N20838 Segment
X20838 N20838 N20839 Segment
X20839 N20839 N20840 Segment
X20840 N20840 N20841 Segment
X20841 N20841 N20842 Segment
X20842 N20842 N20843 Segment
X20843 N20843 N20844 Segment
X20844 N20844 N20845 Segment
X20845 N20845 N20846 Segment
X20846 N20846 N20847 Segment
X20847 N20847 N20848 Segment
X20848 N20848 N20849 Segment
X20849 N20849 N20850 Segment
X20850 N20850 N20851 Segment
X20851 N20851 N20852 Segment
X20852 N20852 N20853 Segment
X20853 N20853 N20854 Segment
X20854 N20854 N20855 Segment
X20855 N20855 N20856 Segment
X20856 N20856 N20857 Segment
X20857 N20857 N20858 Segment
X20858 N20858 N20859 Segment
X20859 N20859 N20860 Segment
X20860 N20860 N20861 Segment
X20861 N20861 N20862 Segment
X20862 N20862 N20863 Segment
X20863 N20863 N20864 Segment
X20864 N20864 N20865 Segment
X20865 N20865 N20866 Segment
X20866 N20866 N20867 Segment
X20867 N20867 N20868 Segment
X20868 N20868 N20869 Segment
X20869 N20869 N20870 Segment
X20870 N20870 N20871 Segment
X20871 N20871 N20872 Segment
X20872 N20872 N20873 Segment
X20873 N20873 N20874 Segment
X20874 N20874 N20875 Segment
X20875 N20875 N20876 Segment
X20876 N20876 N20877 Segment
X20877 N20877 N20878 Segment
X20878 N20878 N20879 Segment
X20879 N20879 N20880 Segment
X20880 N20880 N20881 Segment
X20881 N20881 N20882 Segment
X20882 N20882 N20883 Segment
X20883 N20883 N20884 Segment
X20884 N20884 N20885 Segment
X20885 N20885 N20886 Segment
X20886 N20886 N20887 Segment
X20887 N20887 N20888 Segment
X20888 N20888 N20889 Segment
X20889 N20889 N20890 Segment
X20890 N20890 N20891 Segment
X20891 N20891 N20892 Segment
X20892 N20892 N20893 Segment
X20893 N20893 N20894 Segment
X20894 N20894 N20895 Segment
X20895 N20895 N20896 Segment
X20896 N20896 N20897 Segment
X20897 N20897 N20898 Segment
X20898 N20898 N20899 Segment
X20899 N20899 N20900 Segment
X20900 N20900 N20901 Segment
X20901 N20901 N20902 Segment
X20902 N20902 N20903 Segment
X20903 N20903 N20904 Segment
X20904 N20904 N20905 Segment
X20905 N20905 N20906 Segment
X20906 N20906 N20907 Segment
X20907 N20907 N20908 Segment
X20908 N20908 N20909 Segment
X20909 N20909 N20910 Segment
X20910 N20910 N20911 Segment
X20911 N20911 N20912 Segment
X20912 N20912 N20913 Segment
X20913 N20913 N20914 Segment
X20914 N20914 N20915 Segment
X20915 N20915 N20916 Segment
X20916 N20916 N20917 Segment
X20917 N20917 N20918 Segment
X20918 N20918 N20919 Segment
X20919 N20919 N20920 Segment
X20920 N20920 N20921 Segment
X20921 N20921 N20922 Segment
X20922 N20922 N20923 Segment
X20923 N20923 N20924 Segment
X20924 N20924 N20925 Segment
X20925 N20925 N20926 Segment
X20926 N20926 N20927 Segment
X20927 N20927 N20928 Segment
X20928 N20928 N20929 Segment
X20929 N20929 N20930 Segment
X20930 N20930 N20931 Segment
X20931 N20931 N20932 Segment
X20932 N20932 N20933 Segment
X20933 N20933 N20934 Segment
X20934 N20934 N20935 Segment
X20935 N20935 N20936 Segment
X20936 N20936 N20937 Segment
X20937 N20937 N20938 Segment
X20938 N20938 N20939 Segment
X20939 N20939 N20940 Segment
X20940 N20940 N20941 Segment
X20941 N20941 N20942 Segment
X20942 N20942 N20943 Segment
X20943 N20943 N20944 Segment
X20944 N20944 N20945 Segment
X20945 N20945 N20946 Segment
X20946 N20946 N20947 Segment
X20947 N20947 N20948 Segment
X20948 N20948 N20949 Segment
X20949 N20949 N20950 Segment
X20950 N20950 N20951 Segment
X20951 N20951 N20952 Segment
X20952 N20952 N20953 Segment
X20953 N20953 N20954 Segment
X20954 N20954 N20955 Segment
X20955 N20955 N20956 Segment
X20956 N20956 N20957 Segment
X20957 N20957 N20958 Segment
X20958 N20958 N20959 Segment
X20959 N20959 N20960 Segment
X20960 N20960 N20961 Segment
X20961 N20961 N20962 Segment
X20962 N20962 N20963 Segment
X20963 N20963 N20964 Segment
X20964 N20964 N20965 Segment
X20965 N20965 N20966 Segment
X20966 N20966 N20967 Segment
X20967 N20967 N20968 Segment
X20968 N20968 N20969 Segment
X20969 N20969 N20970 Segment
X20970 N20970 N20971 Segment
X20971 N20971 N20972 Segment
X20972 N20972 N20973 Segment
X20973 N20973 N20974 Segment
X20974 N20974 N20975 Segment
X20975 N20975 N20976 Segment
X20976 N20976 N20977 Segment
X20977 N20977 N20978 Segment
X20978 N20978 N20979 Segment
X20979 N20979 N20980 Segment
X20980 N20980 N20981 Segment
X20981 N20981 N20982 Segment
X20982 N20982 N20983 Segment
X20983 N20983 N20984 Segment
X20984 N20984 N20985 Segment
X20985 N20985 N20986 Segment
X20986 N20986 N20987 Segment
X20987 N20987 N20988 Segment
X20988 N20988 N20989 Segment
X20989 N20989 N20990 Segment
X20990 N20990 N20991 Segment
X20991 N20991 N20992 Segment
X20992 N20992 N20993 Segment
X20993 N20993 N20994 Segment
X20994 N20994 N20995 Segment
X20995 N20995 N20996 Segment
X20996 N20996 N20997 Segment
X20997 N20997 N20998 Segment
X20998 N20998 N20999 Segment
X20999 N20999 N21000 Segment
X21000 N21000 N21001 Segment
X21001 N21001 N21002 Segment
X21002 N21002 N21003 Segment
X21003 N21003 N21004 Segment
X21004 N21004 N21005 Segment
X21005 N21005 N21006 Segment
X21006 N21006 N21007 Segment
X21007 N21007 N21008 Segment
X21008 N21008 N21009 Segment
X21009 N21009 N21010 Segment
X21010 N21010 N21011 Segment
X21011 N21011 N21012 Segment
X21012 N21012 N21013 Segment
X21013 N21013 N21014 Segment
X21014 N21014 N21015 Segment
X21015 N21015 N21016 Segment
X21016 N21016 N21017 Segment
X21017 N21017 N21018 Segment
X21018 N21018 N21019 Segment
X21019 N21019 N21020 Segment
X21020 N21020 N21021 Segment
X21021 N21021 N21022 Segment
X21022 N21022 N21023 Segment
X21023 N21023 N21024 Segment
X21024 N21024 N21025 Segment
X21025 N21025 N21026 Segment
X21026 N21026 N21027 Segment
X21027 N21027 N21028 Segment
X21028 N21028 N21029 Segment
X21029 N21029 N21030 Segment
X21030 N21030 N21031 Segment
X21031 N21031 N21032 Segment
X21032 N21032 N21033 Segment
X21033 N21033 N21034 Segment
X21034 N21034 N21035 Segment
X21035 N21035 N21036 Segment
X21036 N21036 N21037 Segment
X21037 N21037 N21038 Segment
X21038 N21038 N21039 Segment
X21039 N21039 N21040 Segment
X21040 N21040 N21041 Segment
X21041 N21041 N21042 Segment
X21042 N21042 N21043 Segment
X21043 N21043 N21044 Segment
X21044 N21044 N21045 Segment
X21045 N21045 N21046 Segment
X21046 N21046 N21047 Segment
X21047 N21047 N21048 Segment
X21048 N21048 N21049 Segment
X21049 N21049 N21050 Segment
X21050 N21050 N21051 Segment
X21051 N21051 N21052 Segment
X21052 N21052 N21053 Segment
X21053 N21053 N21054 Segment
X21054 N21054 N21055 Segment
X21055 N21055 N21056 Segment
X21056 N21056 N21057 Segment
X21057 N21057 N21058 Segment
X21058 N21058 N21059 Segment
X21059 N21059 N21060 Segment
X21060 N21060 N21061 Segment
X21061 N21061 N21062 Segment
X21062 N21062 N21063 Segment
X21063 N21063 N21064 Segment
X21064 N21064 N21065 Segment
X21065 N21065 N21066 Segment
X21066 N21066 N21067 Segment
X21067 N21067 N21068 Segment
X21068 N21068 N21069 Segment
X21069 N21069 N21070 Segment
X21070 N21070 N21071 Segment
X21071 N21071 N21072 Segment
X21072 N21072 N21073 Segment
X21073 N21073 N21074 Segment
X21074 N21074 N21075 Segment
X21075 N21075 N21076 Segment
X21076 N21076 N21077 Segment
X21077 N21077 N21078 Segment
X21078 N21078 N21079 Segment
X21079 N21079 N21080 Segment
X21080 N21080 N21081 Segment
X21081 N21081 N21082 Segment
X21082 N21082 N21083 Segment
X21083 N21083 N21084 Segment
X21084 N21084 N21085 Segment
X21085 N21085 N21086 Segment
X21086 N21086 N21087 Segment
X21087 N21087 N21088 Segment
X21088 N21088 N21089 Segment
X21089 N21089 N21090 Segment
X21090 N21090 N21091 Segment
X21091 N21091 N21092 Segment
X21092 N21092 N21093 Segment
X21093 N21093 N21094 Segment
X21094 N21094 N21095 Segment
X21095 N21095 N21096 Segment
X21096 N21096 N21097 Segment
X21097 N21097 N21098 Segment
X21098 N21098 N21099 Segment
X21099 N21099 N21100 Segment
X21100 N21100 N21101 Segment
X21101 N21101 N21102 Segment
X21102 N21102 N21103 Segment
X21103 N21103 N21104 Segment
X21104 N21104 N21105 Segment
X21105 N21105 N21106 Segment
X21106 N21106 N21107 Segment
X21107 N21107 N21108 Segment
X21108 N21108 N21109 Segment
X21109 N21109 N21110 Segment
X21110 N21110 N21111 Segment
X21111 N21111 N21112 Segment
X21112 N21112 N21113 Segment
X21113 N21113 N21114 Segment
X21114 N21114 N21115 Segment
X21115 N21115 N21116 Segment
X21116 N21116 N21117 Segment
X21117 N21117 N21118 Segment
X21118 N21118 N21119 Segment
X21119 N21119 N21120 Segment
X21120 N21120 N21121 Segment
X21121 N21121 N21122 Segment
X21122 N21122 N21123 Segment
X21123 N21123 N21124 Segment
X21124 N21124 N21125 Segment
X21125 N21125 N21126 Segment
X21126 N21126 N21127 Segment
X21127 N21127 N21128 Segment
X21128 N21128 N21129 Segment
X21129 N21129 N21130 Segment
X21130 N21130 N21131 Segment
X21131 N21131 N21132 Segment
X21132 N21132 N21133 Segment
X21133 N21133 N21134 Segment
X21134 N21134 N21135 Segment
X21135 N21135 N21136 Segment
X21136 N21136 N21137 Segment
X21137 N21137 N21138 Segment
X21138 N21138 N21139 Segment
X21139 N21139 N21140 Segment
X21140 N21140 N21141 Segment
X21141 N21141 N21142 Segment
X21142 N21142 N21143 Segment
X21143 N21143 N21144 Segment
X21144 N21144 N21145 Segment
X21145 N21145 N21146 Segment
X21146 N21146 N21147 Segment
X21147 N21147 N21148 Segment
X21148 N21148 N21149 Segment
X21149 N21149 N21150 Segment
X21150 N21150 N21151 Segment
X21151 N21151 N21152 Segment
X21152 N21152 N21153 Segment
X21153 N21153 N21154 Segment
X21154 N21154 N21155 Segment
X21155 N21155 N21156 Segment
X21156 N21156 N21157 Segment
X21157 N21157 N21158 Segment
X21158 N21158 N21159 Segment
X21159 N21159 N21160 Segment
X21160 N21160 N21161 Segment
X21161 N21161 N21162 Segment
X21162 N21162 N21163 Segment
X21163 N21163 N21164 Segment
X21164 N21164 N21165 Segment
X21165 N21165 N21166 Segment
X21166 N21166 N21167 Segment
X21167 N21167 N21168 Segment
X21168 N21168 N21169 Segment
X21169 N21169 N21170 Segment
X21170 N21170 N21171 Segment
X21171 N21171 N21172 Segment
X21172 N21172 N21173 Segment
X21173 N21173 N21174 Segment
X21174 N21174 N21175 Segment
X21175 N21175 N21176 Segment
X21176 N21176 N21177 Segment
X21177 N21177 N21178 Segment
X21178 N21178 N21179 Segment
X21179 N21179 N21180 Segment
X21180 N21180 N21181 Segment
X21181 N21181 N21182 Segment
X21182 N21182 N21183 Segment
X21183 N21183 N21184 Segment
X21184 N21184 N21185 Segment
X21185 N21185 N21186 Segment
X21186 N21186 N21187 Segment
X21187 N21187 N21188 Segment
X21188 N21188 N21189 Segment
X21189 N21189 N21190 Segment
X21190 N21190 N21191 Segment
X21191 N21191 N21192 Segment
X21192 N21192 N21193 Segment
X21193 N21193 N21194 Segment
X21194 N21194 N21195 Segment
X21195 N21195 N21196 Segment
X21196 N21196 N21197 Segment
X21197 N21197 N21198 Segment
X21198 N21198 N21199 Segment
X21199 N21199 N21200 Segment
X21200 N21200 N21201 Segment
X21201 N21201 N21202 Segment
X21202 N21202 N21203 Segment
X21203 N21203 N21204 Segment
X21204 N21204 N21205 Segment
X21205 N21205 N21206 Segment
X21206 N21206 N21207 Segment
X21207 N21207 N21208 Segment
X21208 N21208 N21209 Segment
X21209 N21209 N21210 Segment
X21210 N21210 N21211 Segment
X21211 N21211 N21212 Segment
X21212 N21212 N21213 Segment
X21213 N21213 N21214 Segment
X21214 N21214 N21215 Segment
X21215 N21215 N21216 Segment
X21216 N21216 N21217 Segment
X21217 N21217 N21218 Segment
X21218 N21218 N21219 Segment
X21219 N21219 N21220 Segment
X21220 N21220 N21221 Segment
X21221 N21221 N21222 Segment
X21222 N21222 N21223 Segment
X21223 N21223 N21224 Segment
X21224 N21224 N21225 Segment
X21225 N21225 N21226 Segment
X21226 N21226 N21227 Segment
X21227 N21227 N21228 Segment
X21228 N21228 N21229 Segment
X21229 N21229 N21230 Segment
X21230 N21230 N21231 Segment
X21231 N21231 N21232 Segment
X21232 N21232 N21233 Segment
X21233 N21233 N21234 Segment
X21234 N21234 N21235 Segment
X21235 N21235 N21236 Segment
X21236 N21236 N21237 Segment
X21237 N21237 N21238 Segment
X21238 N21238 N21239 Segment
X21239 N21239 N21240 Segment
X21240 N21240 N21241 Segment
X21241 N21241 N21242 Segment
X21242 N21242 N21243 Segment
X21243 N21243 N21244 Segment
X21244 N21244 N21245 Segment
X21245 N21245 N21246 Segment
X21246 N21246 N21247 Segment
X21247 N21247 N21248 Segment
X21248 N21248 N21249 Segment
X21249 N21249 N21250 Segment
X21250 N21250 N21251 Segment
X21251 N21251 N21252 Segment
X21252 N21252 N21253 Segment
X21253 N21253 N21254 Segment
X21254 N21254 N21255 Segment
X21255 N21255 N21256 Segment
X21256 N21256 N21257 Segment
X21257 N21257 N21258 Segment
X21258 N21258 N21259 Segment
X21259 N21259 N21260 Segment
X21260 N21260 N21261 Segment
X21261 N21261 N21262 Segment
X21262 N21262 N21263 Segment
X21263 N21263 N21264 Segment
X21264 N21264 N21265 Segment
X21265 N21265 N21266 Segment
X21266 N21266 N21267 Segment
X21267 N21267 N21268 Segment
X21268 N21268 N21269 Segment
X21269 N21269 N21270 Segment
X21270 N21270 N21271 Segment
X21271 N21271 N21272 Segment
X21272 N21272 N21273 Segment
X21273 N21273 N21274 Segment
X21274 N21274 N21275 Segment
X21275 N21275 N21276 Segment
X21276 N21276 N21277 Segment
X21277 N21277 N21278 Segment
X21278 N21278 N21279 Segment
X21279 N21279 N21280 Segment
X21280 N21280 N21281 Segment
X21281 N21281 N21282 Segment
X21282 N21282 N21283 Segment
X21283 N21283 N21284 Segment
X21284 N21284 N21285 Segment
X21285 N21285 N21286 Segment
X21286 N21286 N21287 Segment
X21287 N21287 N21288 Segment
X21288 N21288 N21289 Segment
X21289 N21289 N21290 Segment
X21290 N21290 N21291 Segment
X21291 N21291 N21292 Segment
X21292 N21292 N21293 Segment
X21293 N21293 N21294 Segment
X21294 N21294 N21295 Segment
X21295 N21295 N21296 Segment
X21296 N21296 N21297 Segment
X21297 N21297 N21298 Segment
X21298 N21298 N21299 Segment
X21299 N21299 N21300 Segment
X21300 N21300 N21301 Segment
X21301 N21301 N21302 Segment
X21302 N21302 N21303 Segment
X21303 N21303 N21304 Segment
X21304 N21304 N21305 Segment
X21305 N21305 N21306 Segment
X21306 N21306 N21307 Segment
X21307 N21307 N21308 Segment
X21308 N21308 N21309 Segment
X21309 N21309 N21310 Segment
X21310 N21310 N21311 Segment
X21311 N21311 N21312 Segment
X21312 N21312 N21313 Segment
X21313 N21313 N21314 Segment
X21314 N21314 N21315 Segment
X21315 N21315 N21316 Segment
X21316 N21316 N21317 Segment
X21317 N21317 N21318 Segment
X21318 N21318 N21319 Segment
X21319 N21319 N21320 Segment
X21320 N21320 N21321 Segment
X21321 N21321 N21322 Segment
X21322 N21322 N21323 Segment
X21323 N21323 N21324 Segment
X21324 N21324 N21325 Segment
X21325 N21325 N21326 Segment
X21326 N21326 N21327 Segment
X21327 N21327 N21328 Segment
X21328 N21328 N21329 Segment
X21329 N21329 N21330 Segment
X21330 N21330 N21331 Segment
X21331 N21331 N21332 Segment
X21332 N21332 N21333 Segment
X21333 N21333 N21334 Segment
X21334 N21334 N21335 Segment
X21335 N21335 N21336 Segment
X21336 N21336 N21337 Segment
X21337 N21337 N21338 Segment
X21338 N21338 N21339 Segment
X21339 N21339 N21340 Segment
X21340 N21340 N21341 Segment
X21341 N21341 N21342 Segment
X21342 N21342 N21343 Segment
X21343 N21343 N21344 Segment
X21344 N21344 N21345 Segment
X21345 N21345 N21346 Segment
X21346 N21346 N21347 Segment
X21347 N21347 N21348 Segment
X21348 N21348 N21349 Segment
X21349 N21349 N21350 Segment
X21350 N21350 N21351 Segment
X21351 N21351 N21352 Segment
X21352 N21352 N21353 Segment
X21353 N21353 N21354 Segment
X21354 N21354 N21355 Segment
X21355 N21355 N21356 Segment
X21356 N21356 N21357 Segment
X21357 N21357 N21358 Segment
X21358 N21358 N21359 Segment
X21359 N21359 N21360 Segment
X21360 N21360 N21361 Segment
X21361 N21361 N21362 Segment
X21362 N21362 N21363 Segment
X21363 N21363 N21364 Segment
X21364 N21364 N21365 Segment
X21365 N21365 N21366 Segment
X21366 N21366 N21367 Segment
X21367 N21367 N21368 Segment
X21368 N21368 N21369 Segment
X21369 N21369 N21370 Segment
X21370 N21370 N21371 Segment
X21371 N21371 N21372 Segment
X21372 N21372 N21373 Segment
X21373 N21373 N21374 Segment
X21374 N21374 N21375 Segment
X21375 N21375 N21376 Segment
X21376 N21376 N21377 Segment
X21377 N21377 N21378 Segment
X21378 N21378 N21379 Segment
X21379 N21379 N21380 Segment
X21380 N21380 N21381 Segment
X21381 N21381 N21382 Segment
X21382 N21382 N21383 Segment
X21383 N21383 N21384 Segment
X21384 N21384 N21385 Segment
X21385 N21385 N21386 Segment
X21386 N21386 N21387 Segment
X21387 N21387 N21388 Segment
X21388 N21388 N21389 Segment
X21389 N21389 N21390 Segment
X21390 N21390 N21391 Segment
X21391 N21391 N21392 Segment
X21392 N21392 N21393 Segment
X21393 N21393 N21394 Segment
X21394 N21394 N21395 Segment
X21395 N21395 N21396 Segment
X21396 N21396 N21397 Segment
X21397 N21397 N21398 Segment
X21398 N21398 N21399 Segment
X21399 N21399 N21400 Segment
X21400 N21400 N21401 Segment
X21401 N21401 N21402 Segment
X21402 N21402 N21403 Segment
X21403 N21403 N21404 Segment
X21404 N21404 N21405 Segment
X21405 N21405 N21406 Segment
X21406 N21406 N21407 Segment
X21407 N21407 N21408 Segment
X21408 N21408 N21409 Segment
X21409 N21409 N21410 Segment
X21410 N21410 N21411 Segment
X21411 N21411 N21412 Segment
X21412 N21412 N21413 Segment
X21413 N21413 N21414 Segment
X21414 N21414 N21415 Segment
X21415 N21415 N21416 Segment
X21416 N21416 N21417 Segment
X21417 N21417 N21418 Segment
X21418 N21418 N21419 Segment
X21419 N21419 N21420 Segment
X21420 N21420 N21421 Segment
X21421 N21421 N21422 Segment
X21422 N21422 N21423 Segment
X21423 N21423 N21424 Segment
X21424 N21424 N21425 Segment
X21425 N21425 N21426 Segment
X21426 N21426 N21427 Segment
X21427 N21427 N21428 Segment
X21428 N21428 N21429 Segment
X21429 N21429 N21430 Segment
X21430 N21430 N21431 Segment
X21431 N21431 N21432 Segment
X21432 N21432 N21433 Segment
X21433 N21433 N21434 Segment
X21434 N21434 N21435 Segment
X21435 N21435 N21436 Segment
X21436 N21436 N21437 Segment
X21437 N21437 N21438 Segment
X21438 N21438 N21439 Segment
X21439 N21439 N21440 Segment
X21440 N21440 N21441 Segment
X21441 N21441 N21442 Segment
X21442 N21442 N21443 Segment
X21443 N21443 N21444 Segment
X21444 N21444 N21445 Segment
X21445 N21445 N21446 Segment
X21446 N21446 N21447 Segment
X21447 N21447 N21448 Segment
X21448 N21448 N21449 Segment
X21449 N21449 N21450 Segment
X21450 N21450 N21451 Segment
X21451 N21451 N21452 Segment
X21452 N21452 N21453 Segment
X21453 N21453 N21454 Segment
X21454 N21454 N21455 Segment
X21455 N21455 N21456 Segment
X21456 N21456 N21457 Segment
X21457 N21457 N21458 Segment
X21458 N21458 N21459 Segment
X21459 N21459 N21460 Segment
X21460 N21460 N21461 Segment
X21461 N21461 N21462 Segment
X21462 N21462 N21463 Segment
X21463 N21463 N21464 Segment
X21464 N21464 N21465 Segment
X21465 N21465 N21466 Segment
X21466 N21466 N21467 Segment
X21467 N21467 N21468 Segment
X21468 N21468 N21469 Segment
X21469 N21469 N21470 Segment
X21470 N21470 N21471 Segment
X21471 N21471 N21472 Segment
X21472 N21472 N21473 Segment
X21473 N21473 N21474 Segment
X21474 N21474 N21475 Segment
X21475 N21475 N21476 Segment
X21476 N21476 N21477 Segment
X21477 N21477 N21478 Segment
X21478 N21478 N21479 Segment
X21479 N21479 N21480 Segment
X21480 N21480 N21481 Segment
X21481 N21481 N21482 Segment
X21482 N21482 N21483 Segment
X21483 N21483 N21484 Segment
X21484 N21484 N21485 Segment
X21485 N21485 N21486 Segment
X21486 N21486 N21487 Segment
X21487 N21487 N21488 Segment
X21488 N21488 N21489 Segment
X21489 N21489 N21490 Segment
X21490 N21490 N21491 Segment
X21491 N21491 N21492 Segment
X21492 N21492 N21493 Segment
X21493 N21493 N21494 Segment
X21494 N21494 N21495 Segment
X21495 N21495 N21496 Segment
X21496 N21496 N21497 Segment
X21497 N21497 N21498 Segment
X21498 N21498 N21499 Segment
X21499 N21499 N21500 Segment
X21500 N21500 N21501 Segment
X21501 N21501 N21502 Segment
X21502 N21502 N21503 Segment
X21503 N21503 N21504 Segment
X21504 N21504 N21505 Segment
X21505 N21505 N21506 Segment
X21506 N21506 N21507 Segment
X21507 N21507 N21508 Segment
X21508 N21508 N21509 Segment
X21509 N21509 N21510 Segment
X21510 N21510 N21511 Segment
X21511 N21511 N21512 Segment
X21512 N21512 N21513 Segment
X21513 N21513 N21514 Segment
X21514 N21514 N21515 Segment
X21515 N21515 N21516 Segment
X21516 N21516 N21517 Segment
X21517 N21517 N21518 Segment
X21518 N21518 N21519 Segment
X21519 N21519 N21520 Segment
X21520 N21520 N21521 Segment
X21521 N21521 N21522 Segment
X21522 N21522 N21523 Segment
X21523 N21523 N21524 Segment
X21524 N21524 N21525 Segment
X21525 N21525 N21526 Segment
X21526 N21526 N21527 Segment
X21527 N21527 N21528 Segment
X21528 N21528 N21529 Segment
X21529 N21529 N21530 Segment
X21530 N21530 N21531 Segment
X21531 N21531 N21532 Segment
X21532 N21532 N21533 Segment
X21533 N21533 N21534 Segment
X21534 N21534 N21535 Segment
X21535 N21535 N21536 Segment
X21536 N21536 N21537 Segment
X21537 N21537 N21538 Segment
X21538 N21538 N21539 Segment
X21539 N21539 N21540 Segment
X21540 N21540 N21541 Segment
X21541 N21541 N21542 Segment
X21542 N21542 N21543 Segment
X21543 N21543 N21544 Segment
X21544 N21544 N21545 Segment
X21545 N21545 N21546 Segment
X21546 N21546 N21547 Segment
X21547 N21547 N21548 Segment
X21548 N21548 N21549 Segment
X21549 N21549 N21550 Segment
X21550 N21550 N21551 Segment
X21551 N21551 N21552 Segment
X21552 N21552 N21553 Segment
X21553 N21553 N21554 Segment
X21554 N21554 N21555 Segment
X21555 N21555 N21556 Segment
X21556 N21556 N21557 Segment
X21557 N21557 N21558 Segment
X21558 N21558 N21559 Segment
X21559 N21559 N21560 Segment
X21560 N21560 N21561 Segment
X21561 N21561 N21562 Segment
X21562 N21562 N21563 Segment
X21563 N21563 N21564 Segment
X21564 N21564 N21565 Segment
X21565 N21565 N21566 Segment
X21566 N21566 N21567 Segment
X21567 N21567 N21568 Segment
X21568 N21568 N21569 Segment
X21569 N21569 N21570 Segment
X21570 N21570 N21571 Segment
X21571 N21571 N21572 Segment
X21572 N21572 N21573 Segment
X21573 N21573 N21574 Segment
X21574 N21574 N21575 Segment
X21575 N21575 N21576 Segment
X21576 N21576 N21577 Segment
X21577 N21577 N21578 Segment
X21578 N21578 N21579 Segment
X21579 N21579 N21580 Segment
X21580 N21580 N21581 Segment
X21581 N21581 N21582 Segment
X21582 N21582 N21583 Segment
X21583 N21583 N21584 Segment
X21584 N21584 N21585 Segment
X21585 N21585 N21586 Segment
X21586 N21586 N21587 Segment
X21587 N21587 N21588 Segment
X21588 N21588 N21589 Segment
X21589 N21589 N21590 Segment
X21590 N21590 N21591 Segment
X21591 N21591 N21592 Segment
X21592 N21592 N21593 Segment
X21593 N21593 N21594 Segment
X21594 N21594 N21595 Segment
X21595 N21595 N21596 Segment
X21596 N21596 N21597 Segment
X21597 N21597 N21598 Segment
X21598 N21598 N21599 Segment
X21599 N21599 N21600 Segment
X21600 N21600 N21601 Segment
X21601 N21601 N21602 Segment
X21602 N21602 N21603 Segment
X21603 N21603 N21604 Segment
X21604 N21604 N21605 Segment
X21605 N21605 N21606 Segment
X21606 N21606 N21607 Segment
X21607 N21607 N21608 Segment
X21608 N21608 N21609 Segment
X21609 N21609 N21610 Segment
X21610 N21610 N21611 Segment
X21611 N21611 N21612 Segment
X21612 N21612 N21613 Segment
X21613 N21613 N21614 Segment
X21614 N21614 N21615 Segment
X21615 N21615 N21616 Segment
X21616 N21616 N21617 Segment
X21617 N21617 N21618 Segment
X21618 N21618 N21619 Segment
X21619 N21619 N21620 Segment
X21620 N21620 N21621 Segment
X21621 N21621 N21622 Segment
X21622 N21622 N21623 Segment
X21623 N21623 N21624 Segment
X21624 N21624 N21625 Segment
X21625 N21625 N21626 Segment
X21626 N21626 N21627 Segment
X21627 N21627 N21628 Segment
X21628 N21628 N21629 Segment
X21629 N21629 N21630 Segment
X21630 N21630 N21631 Segment
X21631 N21631 N21632 Segment
X21632 N21632 N21633 Segment
X21633 N21633 N21634 Segment
X21634 N21634 N21635 Segment
X21635 N21635 N21636 Segment
X21636 N21636 N21637 Segment
X21637 N21637 N21638 Segment
X21638 N21638 N21639 Segment
X21639 N21639 N21640 Segment
X21640 N21640 N21641 Segment
X21641 N21641 N21642 Segment
X21642 N21642 N21643 Segment
X21643 N21643 N21644 Segment
X21644 N21644 N21645 Segment
X21645 N21645 N21646 Segment
X21646 N21646 N21647 Segment
X21647 N21647 N21648 Segment
X21648 N21648 N21649 Segment
X21649 N21649 N21650 Segment
X21650 N21650 N21651 Segment
X21651 N21651 N21652 Segment
X21652 N21652 N21653 Segment
X21653 N21653 N21654 Segment
X21654 N21654 N21655 Segment
X21655 N21655 N21656 Segment
X21656 N21656 N21657 Segment
X21657 N21657 N21658 Segment
X21658 N21658 N21659 Segment
X21659 N21659 N21660 Segment
X21660 N21660 N21661 Segment
X21661 N21661 N21662 Segment
X21662 N21662 N21663 Segment
X21663 N21663 N21664 Segment
X21664 N21664 N21665 Segment
X21665 N21665 N21666 Segment
X21666 N21666 N21667 Segment
X21667 N21667 N21668 Segment
X21668 N21668 N21669 Segment
X21669 N21669 N21670 Segment
X21670 N21670 N21671 Segment
X21671 N21671 N21672 Segment
X21672 N21672 N21673 Segment
X21673 N21673 N21674 Segment
X21674 N21674 N21675 Segment
X21675 N21675 N21676 Segment
X21676 N21676 N21677 Segment
X21677 N21677 N21678 Segment
X21678 N21678 N21679 Segment
X21679 N21679 N21680 Segment
X21680 N21680 N21681 Segment
X21681 N21681 N21682 Segment
X21682 N21682 N21683 Segment
X21683 N21683 N21684 Segment
X21684 N21684 N21685 Segment
X21685 N21685 N21686 Segment
X21686 N21686 N21687 Segment
X21687 N21687 N21688 Segment
X21688 N21688 N21689 Segment
X21689 N21689 N21690 Segment
X21690 N21690 N21691 Segment
X21691 N21691 N21692 Segment
X21692 N21692 N21693 Segment
X21693 N21693 N21694 Segment
X21694 N21694 N21695 Segment
X21695 N21695 N21696 Segment
X21696 N21696 N21697 Segment
X21697 N21697 N21698 Segment
X21698 N21698 N21699 Segment
X21699 N21699 N21700 Segment
X21700 N21700 N21701 Segment
X21701 N21701 N21702 Segment
X21702 N21702 N21703 Segment
X21703 N21703 N21704 Segment
X21704 N21704 N21705 Segment
X21705 N21705 N21706 Segment
X21706 N21706 N21707 Segment
X21707 N21707 N21708 Segment
X21708 N21708 N21709 Segment
X21709 N21709 N21710 Segment
X21710 N21710 N21711 Segment
X21711 N21711 N21712 Segment
X21712 N21712 N21713 Segment
X21713 N21713 N21714 Segment
X21714 N21714 N21715 Segment
X21715 N21715 N21716 Segment
X21716 N21716 N21717 Segment
X21717 N21717 N21718 Segment
X21718 N21718 N21719 Segment
X21719 N21719 N21720 Segment
X21720 N21720 N21721 Segment
X21721 N21721 N21722 Segment
X21722 N21722 N21723 Segment
X21723 N21723 N21724 Segment
X21724 N21724 N21725 Segment
X21725 N21725 N21726 Segment
X21726 N21726 N21727 Segment
X21727 N21727 N21728 Segment
X21728 N21728 N21729 Segment
X21729 N21729 N21730 Segment
X21730 N21730 N21731 Segment
X21731 N21731 N21732 Segment
X21732 N21732 N21733 Segment
X21733 N21733 N21734 Segment
X21734 N21734 N21735 Segment
X21735 N21735 N21736 Segment
X21736 N21736 N21737 Segment
X21737 N21737 N21738 Segment
X21738 N21738 N21739 Segment
X21739 N21739 N21740 Segment
X21740 N21740 N21741 Segment
X21741 N21741 N21742 Segment
X21742 N21742 N21743 Segment
X21743 N21743 N21744 Segment
X21744 N21744 N21745 Segment
X21745 N21745 N21746 Segment
X21746 N21746 N21747 Segment
X21747 N21747 N21748 Segment
X21748 N21748 N21749 Segment
X21749 N21749 N21750 Segment
X21750 N21750 N21751 Segment
X21751 N21751 N21752 Segment
X21752 N21752 N21753 Segment
X21753 N21753 N21754 Segment
X21754 N21754 N21755 Segment
X21755 N21755 N21756 Segment
X21756 N21756 N21757 Segment
X21757 N21757 N21758 Segment
X21758 N21758 N21759 Segment
X21759 N21759 N21760 Segment
X21760 N21760 N21761 Segment
X21761 N21761 N21762 Segment
X21762 N21762 N21763 Segment
X21763 N21763 N21764 Segment
X21764 N21764 N21765 Segment
X21765 N21765 N21766 Segment
X21766 N21766 N21767 Segment
X21767 N21767 N21768 Segment
X21768 N21768 N21769 Segment
X21769 N21769 N21770 Segment
X21770 N21770 N21771 Segment
X21771 N21771 N21772 Segment
X21772 N21772 N21773 Segment
X21773 N21773 N21774 Segment
X21774 N21774 N21775 Segment
X21775 N21775 N21776 Segment
X21776 N21776 N21777 Segment
X21777 N21777 N21778 Segment
X21778 N21778 N21779 Segment
X21779 N21779 N21780 Segment
X21780 N21780 N21781 Segment
X21781 N21781 N21782 Segment
X21782 N21782 N21783 Segment
X21783 N21783 N21784 Segment
X21784 N21784 N21785 Segment
X21785 N21785 N21786 Segment
X21786 N21786 N21787 Segment
X21787 N21787 N21788 Segment
X21788 N21788 N21789 Segment
X21789 N21789 N21790 Segment
X21790 N21790 N21791 Segment
X21791 N21791 N21792 Segment
X21792 N21792 N21793 Segment
X21793 N21793 N21794 Segment
X21794 N21794 N21795 Segment
X21795 N21795 N21796 Segment
X21796 N21796 N21797 Segment
X21797 N21797 N21798 Segment
X21798 N21798 N21799 Segment
X21799 N21799 N21800 Segment
X21800 N21800 N21801 Segment
X21801 N21801 N21802 Segment
X21802 N21802 N21803 Segment
X21803 N21803 N21804 Segment
X21804 N21804 N21805 Segment
X21805 N21805 N21806 Segment
X21806 N21806 N21807 Segment
X21807 N21807 N21808 Segment
X21808 N21808 N21809 Segment
X21809 N21809 N21810 Segment
X21810 N21810 N21811 Segment
X21811 N21811 N21812 Segment
X21812 N21812 N21813 Segment
X21813 N21813 N21814 Segment
X21814 N21814 N21815 Segment
X21815 N21815 N21816 Segment
X21816 N21816 N21817 Segment
X21817 N21817 N21818 Segment
X21818 N21818 N21819 Segment
X21819 N21819 N21820 Segment
X21820 N21820 N21821 Segment
X21821 N21821 N21822 Segment
X21822 N21822 N21823 Segment
X21823 N21823 N21824 Segment
X21824 N21824 N21825 Segment
X21825 N21825 N21826 Segment
X21826 N21826 N21827 Segment
X21827 N21827 N21828 Segment
X21828 N21828 N21829 Segment
X21829 N21829 N21830 Segment
X21830 N21830 N21831 Segment
X21831 N21831 N21832 Segment
X21832 N21832 N21833 Segment
X21833 N21833 N21834 Segment
X21834 N21834 N21835 Segment
X21835 N21835 N21836 Segment
X21836 N21836 N21837 Segment
X21837 N21837 N21838 Segment
X21838 N21838 N21839 Segment
X21839 N21839 N21840 Segment
X21840 N21840 N21841 Segment
X21841 N21841 N21842 Segment
X21842 N21842 N21843 Segment
X21843 N21843 N21844 Segment
X21844 N21844 N21845 Segment
X21845 N21845 N21846 Segment
X21846 N21846 N21847 Segment
X21847 N21847 N21848 Segment
X21848 N21848 N21849 Segment
X21849 N21849 N21850 Segment
X21850 N21850 N21851 Segment
X21851 N21851 N21852 Segment
X21852 N21852 N21853 Segment
X21853 N21853 N21854 Segment
X21854 N21854 N21855 Segment
X21855 N21855 N21856 Segment
X21856 N21856 N21857 Segment
X21857 N21857 N21858 Segment
X21858 N21858 N21859 Segment
X21859 N21859 N21860 Segment
X21860 N21860 N21861 Segment
X21861 N21861 N21862 Segment
X21862 N21862 N21863 Segment
X21863 N21863 N21864 Segment
X21864 N21864 N21865 Segment
X21865 N21865 N21866 Segment
X21866 N21866 N21867 Segment
X21867 N21867 N21868 Segment
X21868 N21868 N21869 Segment
X21869 N21869 N21870 Segment
X21870 N21870 N21871 Segment
X21871 N21871 N21872 Segment
X21872 N21872 N21873 Segment
X21873 N21873 N21874 Segment
X21874 N21874 N21875 Segment
X21875 N21875 N21876 Segment
X21876 N21876 N21877 Segment
X21877 N21877 N21878 Segment
X21878 N21878 N21879 Segment
X21879 N21879 N21880 Segment
X21880 N21880 N21881 Segment
X21881 N21881 N21882 Segment
X21882 N21882 N21883 Segment
X21883 N21883 N21884 Segment
X21884 N21884 N21885 Segment
X21885 N21885 N21886 Segment
X21886 N21886 N21887 Segment
X21887 N21887 N21888 Segment
X21888 N21888 N21889 Segment
X21889 N21889 N21890 Segment
X21890 N21890 N21891 Segment
X21891 N21891 N21892 Segment
X21892 N21892 N21893 Segment
X21893 N21893 N21894 Segment
X21894 N21894 N21895 Segment
X21895 N21895 N21896 Segment
X21896 N21896 N21897 Segment
X21897 N21897 N21898 Segment
X21898 N21898 N21899 Segment
X21899 N21899 N21900 Segment
X21900 N21900 N21901 Segment
X21901 N21901 N21902 Segment
X21902 N21902 N21903 Segment
X21903 N21903 N21904 Segment
X21904 N21904 N21905 Segment
X21905 N21905 N21906 Segment
X21906 N21906 N21907 Segment
X21907 N21907 N21908 Segment
X21908 N21908 N21909 Segment
X21909 N21909 N21910 Segment
X21910 N21910 N21911 Segment
X21911 N21911 N21912 Segment
X21912 N21912 N21913 Segment
X21913 N21913 N21914 Segment
X21914 N21914 N21915 Segment
X21915 N21915 N21916 Segment
X21916 N21916 N21917 Segment
X21917 N21917 N21918 Segment
X21918 N21918 N21919 Segment
X21919 N21919 N21920 Segment
X21920 N21920 N21921 Segment
X21921 N21921 N21922 Segment
X21922 N21922 N21923 Segment
X21923 N21923 N21924 Segment
X21924 N21924 N21925 Segment
X21925 N21925 N21926 Segment
X21926 N21926 N21927 Segment
X21927 N21927 N21928 Segment
X21928 N21928 N21929 Segment
X21929 N21929 N21930 Segment
X21930 N21930 N21931 Segment
X21931 N21931 N21932 Segment
X21932 N21932 N21933 Segment
X21933 N21933 N21934 Segment
X21934 N21934 N21935 Segment
X21935 N21935 N21936 Segment
X21936 N21936 N21937 Segment
X21937 N21937 N21938 Segment
X21938 N21938 N21939 Segment
X21939 N21939 N21940 Segment
X21940 N21940 N21941 Segment
X21941 N21941 N21942 Segment
X21942 N21942 N21943 Segment
X21943 N21943 N21944 Segment
X21944 N21944 N21945 Segment
X21945 N21945 N21946 Segment
X21946 N21946 N21947 Segment
X21947 N21947 N21948 Segment
X21948 N21948 N21949 Segment
X21949 N21949 N21950 Segment
X21950 N21950 N21951 Segment
X21951 N21951 N21952 Segment
X21952 N21952 N21953 Segment
X21953 N21953 N21954 Segment
X21954 N21954 N21955 Segment
X21955 N21955 N21956 Segment
X21956 N21956 N21957 Segment
X21957 N21957 N21958 Segment
X21958 N21958 N21959 Segment
X21959 N21959 N21960 Segment
X21960 N21960 N21961 Segment
X21961 N21961 N21962 Segment
X21962 N21962 N21963 Segment
X21963 N21963 N21964 Segment
X21964 N21964 N21965 Segment
X21965 N21965 N21966 Segment
X21966 N21966 N21967 Segment
X21967 N21967 N21968 Segment
X21968 N21968 N21969 Segment
X21969 N21969 N21970 Segment
X21970 N21970 N21971 Segment
X21971 N21971 N21972 Segment
X21972 N21972 N21973 Segment
X21973 N21973 N21974 Segment
X21974 N21974 N21975 Segment
X21975 N21975 N21976 Segment
X21976 N21976 N21977 Segment
X21977 N21977 N21978 Segment
X21978 N21978 N21979 Segment
X21979 N21979 N21980 Segment
X21980 N21980 N21981 Segment
X21981 N21981 N21982 Segment
X21982 N21982 N21983 Segment
X21983 N21983 N21984 Segment
X21984 N21984 N21985 Segment
X21985 N21985 N21986 Segment
X21986 N21986 N21987 Segment
X21987 N21987 N21988 Segment
X21988 N21988 N21989 Segment
X21989 N21989 N21990 Segment
X21990 N21990 N21991 Segment
X21991 N21991 N21992 Segment
X21992 N21992 N21993 Segment
X21993 N21993 N21994 Segment
X21994 N21994 N21995 Segment
X21995 N21995 N21996 Segment
X21996 N21996 N21997 Segment
X21997 N21997 N21998 Segment
X21998 N21998 N21999 Segment
X21999 N21999 N22000 Segment
X22000 N22000 N22001 Segment
X22001 N22001 N22002 Segment
X22002 N22002 N22003 Segment
X22003 N22003 N22004 Segment
X22004 N22004 N22005 Segment
X22005 N22005 N22006 Segment
X22006 N22006 N22007 Segment
X22007 N22007 N22008 Segment
X22008 N22008 N22009 Segment
X22009 N22009 N22010 Segment
X22010 N22010 N22011 Segment
X22011 N22011 N22012 Segment
X22012 N22012 N22013 Segment
X22013 N22013 N22014 Segment
X22014 N22014 N22015 Segment
X22015 N22015 N22016 Segment
X22016 N22016 N22017 Segment
X22017 N22017 N22018 Segment
X22018 N22018 N22019 Segment
X22019 N22019 N22020 Segment
X22020 N22020 N22021 Segment
X22021 N22021 N22022 Segment
X22022 N22022 N22023 Segment
X22023 N22023 N22024 Segment
X22024 N22024 N22025 Segment
X22025 N22025 N22026 Segment
X22026 N22026 N22027 Segment
X22027 N22027 N22028 Segment
X22028 N22028 N22029 Segment
X22029 N22029 N22030 Segment
X22030 N22030 N22031 Segment
X22031 N22031 N22032 Segment
X22032 N22032 N22033 Segment
X22033 N22033 N22034 Segment
X22034 N22034 N22035 Segment
X22035 N22035 N22036 Segment
X22036 N22036 N22037 Segment
X22037 N22037 N22038 Segment
X22038 N22038 N22039 Segment
X22039 N22039 N22040 Segment
X22040 N22040 N22041 Segment
X22041 N22041 N22042 Segment
X22042 N22042 N22043 Segment
X22043 N22043 N22044 Segment
X22044 N22044 N22045 Segment
X22045 N22045 N22046 Segment
X22046 N22046 N22047 Segment
X22047 N22047 N22048 Segment
X22048 N22048 N22049 Segment
X22049 N22049 N22050 Segment
X22050 N22050 N22051 Segment
X22051 N22051 N22052 Segment
X22052 N22052 N22053 Segment
X22053 N22053 N22054 Segment
X22054 N22054 N22055 Segment
X22055 N22055 N22056 Segment
X22056 N22056 N22057 Segment
X22057 N22057 N22058 Segment
X22058 N22058 N22059 Segment
X22059 N22059 N22060 Segment
X22060 N22060 N22061 Segment
X22061 N22061 N22062 Segment
X22062 N22062 N22063 Segment
X22063 N22063 N22064 Segment
X22064 N22064 N22065 Segment
X22065 N22065 N22066 Segment
X22066 N22066 N22067 Segment
X22067 N22067 N22068 Segment
X22068 N22068 N22069 Segment
X22069 N22069 N22070 Segment
X22070 N22070 N22071 Segment
X22071 N22071 N22072 Segment
X22072 N22072 N22073 Segment
X22073 N22073 N22074 Segment
X22074 N22074 N22075 Segment
X22075 N22075 N22076 Segment
X22076 N22076 N22077 Segment
X22077 N22077 N22078 Segment
X22078 N22078 N22079 Segment
X22079 N22079 N22080 Segment
X22080 N22080 N22081 Segment
X22081 N22081 N22082 Segment
X22082 N22082 N22083 Segment
X22083 N22083 N22084 Segment
X22084 N22084 N22085 Segment
X22085 N22085 N22086 Segment
X22086 N22086 N22087 Segment
X22087 N22087 N22088 Segment
X22088 N22088 N22089 Segment
X22089 N22089 N22090 Segment
X22090 N22090 N22091 Segment
X22091 N22091 N22092 Segment
X22092 N22092 N22093 Segment
X22093 N22093 N22094 Segment
X22094 N22094 N22095 Segment
X22095 N22095 N22096 Segment
X22096 N22096 N22097 Segment
X22097 N22097 N22098 Segment
X22098 N22098 N22099 Segment
X22099 N22099 N22100 Segment
X22100 N22100 N22101 Segment
X22101 N22101 N22102 Segment
X22102 N22102 N22103 Segment
X22103 N22103 N22104 Segment
X22104 N22104 N22105 Segment
X22105 N22105 N22106 Segment
X22106 N22106 N22107 Segment
X22107 N22107 N22108 Segment
X22108 N22108 N22109 Segment
X22109 N22109 N22110 Segment
X22110 N22110 N22111 Segment
X22111 N22111 N22112 Segment
X22112 N22112 N22113 Segment
X22113 N22113 N22114 Segment
X22114 N22114 N22115 Segment
X22115 N22115 N22116 Segment
X22116 N22116 N22117 Segment
X22117 N22117 N22118 Segment
X22118 N22118 N22119 Segment
X22119 N22119 N22120 Segment
X22120 N22120 N22121 Segment
X22121 N22121 N22122 Segment
X22122 N22122 N22123 Segment
X22123 N22123 N22124 Segment
X22124 N22124 N22125 Segment
X22125 N22125 N22126 Segment
X22126 N22126 N22127 Segment
X22127 N22127 N22128 Segment
X22128 N22128 N22129 Segment
X22129 N22129 N22130 Segment
X22130 N22130 N22131 Segment
X22131 N22131 N22132 Segment
X22132 N22132 N22133 Segment
X22133 N22133 N22134 Segment
X22134 N22134 N22135 Segment
X22135 N22135 N22136 Segment
X22136 N22136 N22137 Segment
X22137 N22137 N22138 Segment
X22138 N22138 N22139 Segment
X22139 N22139 N22140 Segment
X22140 N22140 N22141 Segment
X22141 N22141 N22142 Segment
X22142 N22142 N22143 Segment
X22143 N22143 N22144 Segment
X22144 N22144 N22145 Segment
X22145 N22145 N22146 Segment
X22146 N22146 N22147 Segment
X22147 N22147 N22148 Segment
X22148 N22148 N22149 Segment
X22149 N22149 N22150 Segment
X22150 N22150 N22151 Segment
X22151 N22151 N22152 Segment
X22152 N22152 N22153 Segment
X22153 N22153 N22154 Segment
X22154 N22154 N22155 Segment
X22155 N22155 N22156 Segment
X22156 N22156 N22157 Segment
X22157 N22157 N22158 Segment
X22158 N22158 N22159 Segment
X22159 N22159 N22160 Segment
X22160 N22160 N22161 Segment
X22161 N22161 N22162 Segment
X22162 N22162 N22163 Segment
X22163 N22163 N22164 Segment
X22164 N22164 N22165 Segment
X22165 N22165 N22166 Segment
X22166 N22166 N22167 Segment
X22167 N22167 N22168 Segment
X22168 N22168 N22169 Segment
X22169 N22169 N22170 Segment
X22170 N22170 N22171 Segment
X22171 N22171 N22172 Segment
X22172 N22172 N22173 Segment
X22173 N22173 N22174 Segment
X22174 N22174 N22175 Segment
X22175 N22175 N22176 Segment
X22176 N22176 N22177 Segment
X22177 N22177 N22178 Segment
X22178 N22178 N22179 Segment
X22179 N22179 N22180 Segment
X22180 N22180 N22181 Segment
X22181 N22181 N22182 Segment
X22182 N22182 N22183 Segment
X22183 N22183 N22184 Segment
X22184 N22184 N22185 Segment
X22185 N22185 N22186 Segment
X22186 N22186 N22187 Segment
X22187 N22187 N22188 Segment
X22188 N22188 N22189 Segment
X22189 N22189 N22190 Segment
X22190 N22190 N22191 Segment
X22191 N22191 N22192 Segment
X22192 N22192 N22193 Segment
X22193 N22193 N22194 Segment
X22194 N22194 N22195 Segment
X22195 N22195 N22196 Segment
X22196 N22196 N22197 Segment
X22197 N22197 N22198 Segment
X22198 N22198 N22199 Segment
X22199 N22199 N22200 Segment
X22200 N22200 N22201 Segment
X22201 N22201 N22202 Segment
X22202 N22202 N22203 Segment
X22203 N22203 N22204 Segment
X22204 N22204 N22205 Segment
X22205 N22205 N22206 Segment
X22206 N22206 N22207 Segment
X22207 N22207 N22208 Segment
X22208 N22208 N22209 Segment
X22209 N22209 N22210 Segment
X22210 N22210 N22211 Segment
X22211 N22211 N22212 Segment
X22212 N22212 N22213 Segment
X22213 N22213 N22214 Segment
X22214 N22214 N22215 Segment
X22215 N22215 N22216 Segment
X22216 N22216 N22217 Segment
X22217 N22217 N22218 Segment
X22218 N22218 N22219 Segment
X22219 N22219 N22220 Segment
X22220 N22220 N22221 Segment
X22221 N22221 N22222 Segment
X22222 N22222 N22223 Segment
X22223 N22223 N22224 Segment
X22224 N22224 N22225 Segment
X22225 N22225 N22226 Segment
X22226 N22226 N22227 Segment
X22227 N22227 N22228 Segment
X22228 N22228 N22229 Segment
X22229 N22229 N22230 Segment
X22230 N22230 N22231 Segment
X22231 N22231 N22232 Segment
X22232 N22232 N22233 Segment
X22233 N22233 N22234 Segment
X22234 N22234 N22235 Segment
X22235 N22235 N22236 Segment
X22236 N22236 N22237 Segment
X22237 N22237 N22238 Segment
X22238 N22238 N22239 Segment
X22239 N22239 N22240 Segment
X22240 N22240 N22241 Segment
X22241 N22241 N22242 Segment
X22242 N22242 N22243 Segment
X22243 N22243 N22244 Segment
X22244 N22244 N22245 Segment
X22245 N22245 N22246 Segment
X22246 N22246 N22247 Segment
X22247 N22247 N22248 Segment
X22248 N22248 N22249 Segment
X22249 N22249 N22250 Segment
X22250 N22250 N22251 Segment
X22251 N22251 N22252 Segment
X22252 N22252 N22253 Segment
X22253 N22253 N22254 Segment
X22254 N22254 N22255 Segment
X22255 N22255 N22256 Segment
X22256 N22256 N22257 Segment
X22257 N22257 N22258 Segment
X22258 N22258 N22259 Segment
X22259 N22259 N22260 Segment
X22260 N22260 N22261 Segment
X22261 N22261 N22262 Segment
X22262 N22262 N22263 Segment
X22263 N22263 N22264 Segment
X22264 N22264 N22265 Segment
X22265 N22265 N22266 Segment
X22266 N22266 N22267 Segment
X22267 N22267 N22268 Segment
X22268 N22268 N22269 Segment
X22269 N22269 N22270 Segment
X22270 N22270 N22271 Segment
X22271 N22271 N22272 Segment
X22272 N22272 N22273 Segment
X22273 N22273 N22274 Segment
X22274 N22274 N22275 Segment
X22275 N22275 N22276 Segment
X22276 N22276 N22277 Segment
X22277 N22277 N22278 Segment
X22278 N22278 N22279 Segment
X22279 N22279 N22280 Segment
X22280 N22280 N22281 Segment
X22281 N22281 N22282 Segment
X22282 N22282 N22283 Segment
X22283 N22283 N22284 Segment
X22284 N22284 N22285 Segment
X22285 N22285 N22286 Segment
X22286 N22286 N22287 Segment
X22287 N22287 N22288 Segment
X22288 N22288 N22289 Segment
X22289 N22289 N22290 Segment
X22290 N22290 N22291 Segment
X22291 N22291 N22292 Segment
X22292 N22292 N22293 Segment
X22293 N22293 N22294 Segment
X22294 N22294 N22295 Segment
X22295 N22295 N22296 Segment
X22296 N22296 N22297 Segment
X22297 N22297 N22298 Segment
X22298 N22298 N22299 Segment
X22299 N22299 N22300 Segment
X22300 N22300 N22301 Segment
X22301 N22301 N22302 Segment
X22302 N22302 N22303 Segment
X22303 N22303 N22304 Segment
X22304 N22304 N22305 Segment
X22305 N22305 N22306 Segment
X22306 N22306 N22307 Segment
X22307 N22307 N22308 Segment
X22308 N22308 N22309 Segment
X22309 N22309 N22310 Segment
X22310 N22310 N22311 Segment
X22311 N22311 N22312 Segment
X22312 N22312 N22313 Segment
X22313 N22313 N22314 Segment
X22314 N22314 N22315 Segment
X22315 N22315 N22316 Segment
X22316 N22316 N22317 Segment
X22317 N22317 N22318 Segment
X22318 N22318 N22319 Segment
X22319 N22319 N22320 Segment
X22320 N22320 N22321 Segment
X22321 N22321 N22322 Segment
X22322 N22322 N22323 Segment
X22323 N22323 N22324 Segment
X22324 N22324 N22325 Segment
X22325 N22325 N22326 Segment
X22326 N22326 N22327 Segment
X22327 N22327 N22328 Segment
X22328 N22328 N22329 Segment
X22329 N22329 N22330 Segment
X22330 N22330 N22331 Segment
X22331 N22331 N22332 Segment
X22332 N22332 N22333 Segment
X22333 N22333 N22334 Segment
X22334 N22334 N22335 Segment
X22335 N22335 N22336 Segment
X22336 N22336 N22337 Segment
X22337 N22337 N22338 Segment
X22338 N22338 N22339 Segment
X22339 N22339 N22340 Segment
X22340 N22340 N22341 Segment
X22341 N22341 N22342 Segment
X22342 N22342 N22343 Segment
X22343 N22343 N22344 Segment
X22344 N22344 N22345 Segment
X22345 N22345 N22346 Segment
X22346 N22346 N22347 Segment
X22347 N22347 N22348 Segment
X22348 N22348 N22349 Segment
X22349 N22349 N22350 Segment
X22350 N22350 N22351 Segment
X22351 N22351 N22352 Segment
X22352 N22352 N22353 Segment
X22353 N22353 N22354 Segment
X22354 N22354 N22355 Segment
X22355 N22355 N22356 Segment
X22356 N22356 N22357 Segment
X22357 N22357 N22358 Segment
X22358 N22358 N22359 Segment
X22359 N22359 N22360 Segment
X22360 N22360 N22361 Segment
X22361 N22361 N22362 Segment
X22362 N22362 N22363 Segment
X22363 N22363 N22364 Segment
X22364 N22364 N22365 Segment
X22365 N22365 N22366 Segment
X22366 N22366 N22367 Segment
X22367 N22367 N22368 Segment
X22368 N22368 N22369 Segment
X22369 N22369 N22370 Segment
X22370 N22370 N22371 Segment
X22371 N22371 N22372 Segment
X22372 N22372 N22373 Segment
X22373 N22373 N22374 Segment
X22374 N22374 N22375 Segment
X22375 N22375 N22376 Segment
X22376 N22376 N22377 Segment
X22377 N22377 N22378 Segment
X22378 N22378 N22379 Segment
X22379 N22379 N22380 Segment
X22380 N22380 N22381 Segment
X22381 N22381 N22382 Segment
X22382 N22382 N22383 Segment
X22383 N22383 N22384 Segment
X22384 N22384 N22385 Segment
X22385 N22385 N22386 Segment
X22386 N22386 N22387 Segment
X22387 N22387 N22388 Segment
X22388 N22388 N22389 Segment
X22389 N22389 N22390 Segment
X22390 N22390 N22391 Segment
X22391 N22391 N22392 Segment
X22392 N22392 N22393 Segment
X22393 N22393 N22394 Segment
X22394 N22394 N22395 Segment
X22395 N22395 N22396 Segment
X22396 N22396 N22397 Segment
X22397 N22397 N22398 Segment
X22398 N22398 N22399 Segment
X22399 N22399 N22400 Segment
X22400 N22400 N22401 Segment
X22401 N22401 N22402 Segment
X22402 N22402 N22403 Segment
X22403 N22403 N22404 Segment
X22404 N22404 N22405 Segment
X22405 N22405 N22406 Segment
X22406 N22406 N22407 Segment
X22407 N22407 N22408 Segment
X22408 N22408 N22409 Segment
X22409 N22409 N22410 Segment
X22410 N22410 N22411 Segment
X22411 N22411 N22412 Segment
X22412 N22412 N22413 Segment
X22413 N22413 N22414 Segment
X22414 N22414 N22415 Segment
X22415 N22415 N22416 Segment
X22416 N22416 N22417 Segment
X22417 N22417 N22418 Segment
X22418 N22418 N22419 Segment
X22419 N22419 N22420 Segment
X22420 N22420 N22421 Segment
X22421 N22421 N22422 Segment
X22422 N22422 N22423 Segment
X22423 N22423 N22424 Segment
X22424 N22424 N22425 Segment
X22425 N22425 N22426 Segment
X22426 N22426 N22427 Segment
X22427 N22427 N22428 Segment
X22428 N22428 N22429 Segment
X22429 N22429 N22430 Segment
X22430 N22430 N22431 Segment
X22431 N22431 N22432 Segment
X22432 N22432 N22433 Segment
X22433 N22433 N22434 Segment
X22434 N22434 N22435 Segment
X22435 N22435 N22436 Segment
X22436 N22436 N22437 Segment
X22437 N22437 N22438 Segment
X22438 N22438 N22439 Segment
X22439 N22439 N22440 Segment
X22440 N22440 N22441 Segment
X22441 N22441 N22442 Segment
X22442 N22442 N22443 Segment
X22443 N22443 N22444 Segment
X22444 N22444 N22445 Segment
X22445 N22445 N22446 Segment
X22446 N22446 N22447 Segment
X22447 N22447 N22448 Segment
X22448 N22448 N22449 Segment
X22449 N22449 N22450 Segment
X22450 N22450 N22451 Segment
X22451 N22451 N22452 Segment
X22452 N22452 N22453 Segment
X22453 N22453 N22454 Segment
X22454 N22454 N22455 Segment
X22455 N22455 N22456 Segment
X22456 N22456 N22457 Segment
X22457 N22457 N22458 Segment
X22458 N22458 N22459 Segment
X22459 N22459 N22460 Segment
X22460 N22460 N22461 Segment
X22461 N22461 N22462 Segment
X22462 N22462 N22463 Segment
X22463 N22463 N22464 Segment
X22464 N22464 N22465 Segment
X22465 N22465 N22466 Segment
X22466 N22466 N22467 Segment
X22467 N22467 N22468 Segment
X22468 N22468 N22469 Segment
X22469 N22469 N22470 Segment
X22470 N22470 N22471 Segment
X22471 N22471 N22472 Segment
X22472 N22472 N22473 Segment
X22473 N22473 N22474 Segment
X22474 N22474 N22475 Segment
X22475 N22475 N22476 Segment
X22476 N22476 N22477 Segment
X22477 N22477 N22478 Segment
X22478 N22478 N22479 Segment
X22479 N22479 N22480 Segment
X22480 N22480 N22481 Segment
X22481 N22481 N22482 Segment
X22482 N22482 N22483 Segment
X22483 N22483 N22484 Segment
X22484 N22484 N22485 Segment
X22485 N22485 N22486 Segment
X22486 N22486 N22487 Segment
X22487 N22487 N22488 Segment
X22488 N22488 N22489 Segment
X22489 N22489 N22490 Segment
X22490 N22490 N22491 Segment
X22491 N22491 N22492 Segment
X22492 N22492 N22493 Segment
X22493 N22493 N22494 Segment
X22494 N22494 N22495 Segment
X22495 N22495 N22496 Segment
X22496 N22496 N22497 Segment
X22497 N22497 N22498 Segment
X22498 N22498 N22499 Segment
X22499 N22499 N22500 Segment
X22500 N22500 N22501 Segment
X22501 N22501 N22502 Segment
X22502 N22502 N22503 Segment
X22503 N22503 N22504 Segment
X22504 N22504 N22505 Segment
X22505 N22505 N22506 Segment
X22506 N22506 N22507 Segment
X22507 N22507 N22508 Segment
X22508 N22508 N22509 Segment
X22509 N22509 N22510 Segment
X22510 N22510 N22511 Segment
X22511 N22511 N22512 Segment
X22512 N22512 N22513 Segment
X22513 N22513 N22514 Segment
X22514 N22514 N22515 Segment
X22515 N22515 N22516 Segment
X22516 N22516 N22517 Segment
X22517 N22517 N22518 Segment
X22518 N22518 N22519 Segment
X22519 N22519 N22520 Segment
X22520 N22520 N22521 Segment
X22521 N22521 N22522 Segment
X22522 N22522 N22523 Segment
X22523 N22523 N22524 Segment
X22524 N22524 N22525 Segment
X22525 N22525 N22526 Segment
X22526 N22526 N22527 Segment
X22527 N22527 N22528 Segment
X22528 N22528 N22529 Segment
X22529 N22529 N22530 Segment
X22530 N22530 N22531 Segment
X22531 N22531 N22532 Segment
X22532 N22532 N22533 Segment
X22533 N22533 N22534 Segment
X22534 N22534 N22535 Segment
X22535 N22535 N22536 Segment
X22536 N22536 N22537 Segment
X22537 N22537 N22538 Segment
X22538 N22538 N22539 Segment
X22539 N22539 N22540 Segment
X22540 N22540 N22541 Segment
X22541 N22541 N22542 Segment
X22542 N22542 N22543 Segment
X22543 N22543 N22544 Segment
X22544 N22544 N22545 Segment
X22545 N22545 N22546 Segment
X22546 N22546 N22547 Segment
X22547 N22547 N22548 Segment
X22548 N22548 N22549 Segment
X22549 N22549 N22550 Segment
X22550 N22550 N22551 Segment
X22551 N22551 N22552 Segment
X22552 N22552 N22553 Segment
X22553 N22553 N22554 Segment
X22554 N22554 N22555 Segment
X22555 N22555 N22556 Segment
X22556 N22556 N22557 Segment
X22557 N22557 N22558 Segment
X22558 N22558 N22559 Segment
X22559 N22559 N22560 Segment
X22560 N22560 N22561 Segment
X22561 N22561 N22562 Segment
X22562 N22562 N22563 Segment
X22563 N22563 N22564 Segment
X22564 N22564 N22565 Segment
X22565 N22565 N22566 Segment
X22566 N22566 N22567 Segment
X22567 N22567 N22568 Segment
X22568 N22568 N22569 Segment
X22569 N22569 N22570 Segment
X22570 N22570 N22571 Segment
X22571 N22571 N22572 Segment
X22572 N22572 N22573 Segment
X22573 N22573 N22574 Segment
X22574 N22574 N22575 Segment
X22575 N22575 N22576 Segment
X22576 N22576 N22577 Segment
X22577 N22577 N22578 Segment
X22578 N22578 N22579 Segment
X22579 N22579 N22580 Segment
X22580 N22580 N22581 Segment
X22581 N22581 N22582 Segment
X22582 N22582 N22583 Segment
X22583 N22583 N22584 Segment
X22584 N22584 N22585 Segment
X22585 N22585 N22586 Segment
X22586 N22586 N22587 Segment
X22587 N22587 N22588 Segment
X22588 N22588 N22589 Segment
X22589 N22589 N22590 Segment
X22590 N22590 N22591 Segment
X22591 N22591 N22592 Segment
X22592 N22592 N22593 Segment
X22593 N22593 N22594 Segment
X22594 N22594 N22595 Segment
X22595 N22595 N22596 Segment
X22596 N22596 N22597 Segment
X22597 N22597 N22598 Segment
X22598 N22598 N22599 Segment
X22599 N22599 N22600 Segment
X22600 N22600 N22601 Segment
X22601 N22601 N22602 Segment
X22602 N22602 N22603 Segment
X22603 N22603 N22604 Segment
X22604 N22604 N22605 Segment
X22605 N22605 N22606 Segment
X22606 N22606 N22607 Segment
X22607 N22607 N22608 Segment
X22608 N22608 N22609 Segment
X22609 N22609 N22610 Segment
X22610 N22610 N22611 Segment
X22611 N22611 N22612 Segment
X22612 N22612 N22613 Segment
X22613 N22613 N22614 Segment
X22614 N22614 N22615 Segment
X22615 N22615 N22616 Segment
X22616 N22616 N22617 Segment
X22617 N22617 N22618 Segment
X22618 N22618 N22619 Segment
X22619 N22619 N22620 Segment
X22620 N22620 N22621 Segment
X22621 N22621 N22622 Segment
X22622 N22622 N22623 Segment
X22623 N22623 N22624 Segment
X22624 N22624 N22625 Segment
X22625 N22625 N22626 Segment
X22626 N22626 N22627 Segment
X22627 N22627 N22628 Segment
X22628 N22628 N22629 Segment
X22629 N22629 N22630 Segment
X22630 N22630 N22631 Segment
X22631 N22631 N22632 Segment
X22632 N22632 N22633 Segment
X22633 N22633 N22634 Segment
X22634 N22634 N22635 Segment
X22635 N22635 N22636 Segment
X22636 N22636 N22637 Segment
X22637 N22637 N22638 Segment
X22638 N22638 N22639 Segment
X22639 N22639 N22640 Segment
X22640 N22640 N22641 Segment
X22641 N22641 N22642 Segment
X22642 N22642 N22643 Segment
X22643 N22643 N22644 Segment
X22644 N22644 N22645 Segment
X22645 N22645 N22646 Segment
X22646 N22646 N22647 Segment
X22647 N22647 N22648 Segment
X22648 N22648 N22649 Segment
X22649 N22649 N22650 Segment
X22650 N22650 N22651 Segment
X22651 N22651 N22652 Segment
X22652 N22652 N22653 Segment
X22653 N22653 N22654 Segment
X22654 N22654 N22655 Segment
X22655 N22655 N22656 Segment
X22656 N22656 N22657 Segment
X22657 N22657 N22658 Segment
X22658 N22658 N22659 Segment
X22659 N22659 N22660 Segment
X22660 N22660 N22661 Segment
X22661 N22661 N22662 Segment
X22662 N22662 N22663 Segment
X22663 N22663 N22664 Segment
X22664 N22664 N22665 Segment
X22665 N22665 N22666 Segment
X22666 N22666 N22667 Segment
X22667 N22667 N22668 Segment
X22668 N22668 N22669 Segment
X22669 N22669 N22670 Segment
X22670 N22670 N22671 Segment
X22671 N22671 N22672 Segment
X22672 N22672 N22673 Segment
X22673 N22673 N22674 Segment
X22674 N22674 N22675 Segment
X22675 N22675 N22676 Segment
X22676 N22676 N22677 Segment
X22677 N22677 N22678 Segment
X22678 N22678 N22679 Segment
X22679 N22679 N22680 Segment
X22680 N22680 N22681 Segment
X22681 N22681 N22682 Segment
X22682 N22682 N22683 Segment
X22683 N22683 N22684 Segment
X22684 N22684 N22685 Segment
X22685 N22685 N22686 Segment
X22686 N22686 N22687 Segment
X22687 N22687 N22688 Segment
X22688 N22688 N22689 Segment
X22689 N22689 N22690 Segment
X22690 N22690 N22691 Segment
X22691 N22691 N22692 Segment
X22692 N22692 N22693 Segment
X22693 N22693 N22694 Segment
X22694 N22694 N22695 Segment
X22695 N22695 N22696 Segment
X22696 N22696 N22697 Segment
X22697 N22697 N22698 Segment
X22698 N22698 N22699 Segment
X22699 N22699 N22700 Segment
X22700 N22700 N22701 Segment
X22701 N22701 N22702 Segment
X22702 N22702 N22703 Segment
X22703 N22703 N22704 Segment
X22704 N22704 N22705 Segment
X22705 N22705 N22706 Segment
X22706 N22706 N22707 Segment
X22707 N22707 N22708 Segment
X22708 N22708 N22709 Segment
X22709 N22709 N22710 Segment
X22710 N22710 N22711 Segment
X22711 N22711 N22712 Segment
X22712 N22712 N22713 Segment
X22713 N22713 N22714 Segment
X22714 N22714 N22715 Segment
X22715 N22715 N22716 Segment
X22716 N22716 N22717 Segment
X22717 N22717 N22718 Segment
X22718 N22718 N22719 Segment
X22719 N22719 N22720 Segment
X22720 N22720 N22721 Segment
X22721 N22721 N22722 Segment
X22722 N22722 N22723 Segment
X22723 N22723 N22724 Segment
X22724 N22724 N22725 Segment
X22725 N22725 N22726 Segment
X22726 N22726 N22727 Segment
X22727 N22727 N22728 Segment
X22728 N22728 N22729 Segment
X22729 N22729 N22730 Segment
X22730 N22730 N22731 Segment
X22731 N22731 N22732 Segment
X22732 N22732 N22733 Segment
X22733 N22733 N22734 Segment
X22734 N22734 N22735 Segment
X22735 N22735 N22736 Segment
X22736 N22736 N22737 Segment
X22737 N22737 N22738 Segment
X22738 N22738 N22739 Segment
X22739 N22739 N22740 Segment
X22740 N22740 N22741 Segment
X22741 N22741 N22742 Segment
X22742 N22742 N22743 Segment
X22743 N22743 N22744 Segment
X22744 N22744 N22745 Segment
X22745 N22745 N22746 Segment
X22746 N22746 N22747 Segment
X22747 N22747 N22748 Segment
X22748 N22748 N22749 Segment
X22749 N22749 N22750 Segment
X22750 N22750 N22751 Segment
X22751 N22751 N22752 Segment
X22752 N22752 N22753 Segment
X22753 N22753 N22754 Segment
X22754 N22754 N22755 Segment
X22755 N22755 N22756 Segment
X22756 N22756 N22757 Segment
X22757 N22757 N22758 Segment
X22758 N22758 N22759 Segment
X22759 N22759 N22760 Segment
X22760 N22760 N22761 Segment
X22761 N22761 N22762 Segment
X22762 N22762 N22763 Segment
X22763 N22763 N22764 Segment
X22764 N22764 N22765 Segment
X22765 N22765 N22766 Segment
X22766 N22766 N22767 Segment
X22767 N22767 N22768 Segment
X22768 N22768 N22769 Segment
X22769 N22769 N22770 Segment
X22770 N22770 N22771 Segment
X22771 N22771 N22772 Segment
X22772 N22772 N22773 Segment
X22773 N22773 N22774 Segment
X22774 N22774 N22775 Segment
X22775 N22775 N22776 Segment
X22776 N22776 N22777 Segment
X22777 N22777 N22778 Segment
X22778 N22778 N22779 Segment
X22779 N22779 N22780 Segment
X22780 N22780 N22781 Segment
X22781 N22781 N22782 Segment
X22782 N22782 N22783 Segment
X22783 N22783 N22784 Segment
X22784 N22784 N22785 Segment
X22785 N22785 N22786 Segment
X22786 N22786 N22787 Segment
X22787 N22787 N22788 Segment
X22788 N22788 N22789 Segment
X22789 N22789 N22790 Segment
X22790 N22790 N22791 Segment
X22791 N22791 N22792 Segment
X22792 N22792 N22793 Segment
X22793 N22793 N22794 Segment
X22794 N22794 N22795 Segment
X22795 N22795 N22796 Segment
X22796 N22796 N22797 Segment
X22797 N22797 N22798 Segment
X22798 N22798 N22799 Segment
X22799 N22799 N22800 Segment
X22800 N22800 N22801 Segment
X22801 N22801 N22802 Segment
X22802 N22802 N22803 Segment
X22803 N22803 N22804 Segment
X22804 N22804 N22805 Segment
X22805 N22805 N22806 Segment
X22806 N22806 N22807 Segment
X22807 N22807 N22808 Segment
X22808 N22808 N22809 Segment
X22809 N22809 N22810 Segment
X22810 N22810 N22811 Segment
X22811 N22811 N22812 Segment
X22812 N22812 N22813 Segment
X22813 N22813 N22814 Segment
X22814 N22814 N22815 Segment
X22815 N22815 N22816 Segment
X22816 N22816 N22817 Segment
X22817 N22817 N22818 Segment
X22818 N22818 N22819 Segment
X22819 N22819 N22820 Segment
X22820 N22820 N22821 Segment
X22821 N22821 N22822 Segment
X22822 N22822 N22823 Segment
X22823 N22823 N22824 Segment
X22824 N22824 N22825 Segment
X22825 N22825 N22826 Segment
X22826 N22826 N22827 Segment
X22827 N22827 N22828 Segment
X22828 N22828 N22829 Segment
X22829 N22829 N22830 Segment
X22830 N22830 N22831 Segment
X22831 N22831 N22832 Segment
X22832 N22832 N22833 Segment
X22833 N22833 N22834 Segment
X22834 N22834 N22835 Segment
X22835 N22835 N22836 Segment
X22836 N22836 N22837 Segment
X22837 N22837 N22838 Segment
X22838 N22838 N22839 Segment
X22839 N22839 N22840 Segment
X22840 N22840 N22841 Segment
X22841 N22841 N22842 Segment
X22842 N22842 N22843 Segment
X22843 N22843 N22844 Segment
X22844 N22844 N22845 Segment
X22845 N22845 N22846 Segment
X22846 N22846 N22847 Segment
X22847 N22847 N22848 Segment
X22848 N22848 N22849 Segment
X22849 N22849 N22850 Segment
X22850 N22850 N22851 Segment
X22851 N22851 N22852 Segment
X22852 N22852 N22853 Segment
X22853 N22853 N22854 Segment
X22854 N22854 N22855 Segment
X22855 N22855 N22856 Segment
X22856 N22856 N22857 Segment
X22857 N22857 N22858 Segment
X22858 N22858 N22859 Segment
X22859 N22859 N22860 Segment
X22860 N22860 N22861 Segment
X22861 N22861 N22862 Segment
X22862 N22862 N22863 Segment
X22863 N22863 N22864 Segment
X22864 N22864 N22865 Segment
X22865 N22865 N22866 Segment
X22866 N22866 N22867 Segment
X22867 N22867 N22868 Segment
X22868 N22868 N22869 Segment
X22869 N22869 N22870 Segment
X22870 N22870 N22871 Segment
X22871 N22871 N22872 Segment
X22872 N22872 N22873 Segment
X22873 N22873 N22874 Segment
X22874 N22874 N22875 Segment
X22875 N22875 N22876 Segment
X22876 N22876 N22877 Segment
X22877 N22877 N22878 Segment
X22878 N22878 N22879 Segment
X22879 N22879 N22880 Segment
X22880 N22880 N22881 Segment
X22881 N22881 N22882 Segment
X22882 N22882 N22883 Segment
X22883 N22883 N22884 Segment
X22884 N22884 N22885 Segment
X22885 N22885 N22886 Segment
X22886 N22886 N22887 Segment
X22887 N22887 N22888 Segment
X22888 N22888 N22889 Segment
X22889 N22889 N22890 Segment
X22890 N22890 N22891 Segment
X22891 N22891 N22892 Segment
X22892 N22892 N22893 Segment
X22893 N22893 N22894 Segment
X22894 N22894 N22895 Segment
X22895 N22895 N22896 Segment
X22896 N22896 N22897 Segment
X22897 N22897 N22898 Segment
X22898 N22898 N22899 Segment
X22899 N22899 N22900 Segment
X22900 N22900 N22901 Segment
X22901 N22901 N22902 Segment
X22902 N22902 N22903 Segment
X22903 N22903 N22904 Segment
X22904 N22904 N22905 Segment
X22905 N22905 N22906 Segment
X22906 N22906 N22907 Segment
X22907 N22907 N22908 Segment
X22908 N22908 N22909 Segment
X22909 N22909 N22910 Segment
X22910 N22910 N22911 Segment
X22911 N22911 N22912 Segment
X22912 N22912 N22913 Segment
X22913 N22913 N22914 Segment
X22914 N22914 N22915 Segment
X22915 N22915 N22916 Segment
X22916 N22916 N22917 Segment
X22917 N22917 N22918 Segment
X22918 N22918 N22919 Segment
X22919 N22919 N22920 Segment
X22920 N22920 N22921 Segment
X22921 N22921 N22922 Segment
X22922 N22922 N22923 Segment
X22923 N22923 N22924 Segment
X22924 N22924 N22925 Segment
X22925 N22925 N22926 Segment
X22926 N22926 N22927 Segment
X22927 N22927 N22928 Segment
X22928 N22928 N22929 Segment
X22929 N22929 N22930 Segment
X22930 N22930 N22931 Segment
X22931 N22931 N22932 Segment
X22932 N22932 N22933 Segment
X22933 N22933 N22934 Segment
X22934 N22934 N22935 Segment
X22935 N22935 N22936 Segment
X22936 N22936 N22937 Segment
X22937 N22937 N22938 Segment
X22938 N22938 N22939 Segment
X22939 N22939 N22940 Segment
X22940 N22940 N22941 Segment
X22941 N22941 N22942 Segment
X22942 N22942 N22943 Segment
X22943 N22943 N22944 Segment
X22944 N22944 N22945 Segment
X22945 N22945 N22946 Segment
X22946 N22946 N22947 Segment
X22947 N22947 N22948 Segment
X22948 N22948 N22949 Segment
X22949 N22949 N22950 Segment
X22950 N22950 N22951 Segment
X22951 N22951 N22952 Segment
X22952 N22952 N22953 Segment
X22953 N22953 N22954 Segment
X22954 N22954 N22955 Segment
X22955 N22955 N22956 Segment
X22956 N22956 N22957 Segment
X22957 N22957 N22958 Segment
X22958 N22958 N22959 Segment
X22959 N22959 N22960 Segment
X22960 N22960 N22961 Segment
X22961 N22961 N22962 Segment
X22962 N22962 N22963 Segment
X22963 N22963 N22964 Segment
X22964 N22964 N22965 Segment
X22965 N22965 N22966 Segment
X22966 N22966 N22967 Segment
X22967 N22967 N22968 Segment
X22968 N22968 N22969 Segment
X22969 N22969 N22970 Segment
X22970 N22970 N22971 Segment
X22971 N22971 N22972 Segment
X22972 N22972 N22973 Segment
X22973 N22973 N22974 Segment
X22974 N22974 N22975 Segment
X22975 N22975 N22976 Segment
X22976 N22976 N22977 Segment
X22977 N22977 N22978 Segment
X22978 N22978 N22979 Segment
X22979 N22979 N22980 Segment
X22980 N22980 N22981 Segment
X22981 N22981 N22982 Segment
X22982 N22982 N22983 Segment
X22983 N22983 N22984 Segment
X22984 N22984 N22985 Segment
X22985 N22985 N22986 Segment
X22986 N22986 N22987 Segment
X22987 N22987 N22988 Segment
X22988 N22988 N22989 Segment
X22989 N22989 N22990 Segment
X22990 N22990 N22991 Segment
X22991 N22991 N22992 Segment
X22992 N22992 N22993 Segment
X22993 N22993 N22994 Segment
X22994 N22994 N22995 Segment
X22995 N22995 N22996 Segment
X22996 N22996 N22997 Segment
X22997 N22997 N22998 Segment
X22998 N22998 N22999 Segment
X22999 N22999 N23000 Segment
X23000 N23000 N23001 Segment
X23001 N23001 N23002 Segment
X23002 N23002 N23003 Segment
X23003 N23003 N23004 Segment
X23004 N23004 N23005 Segment
X23005 N23005 N23006 Segment
X23006 N23006 N23007 Segment
X23007 N23007 N23008 Segment
X23008 N23008 N23009 Segment
X23009 N23009 N23010 Segment
X23010 N23010 N23011 Segment
X23011 N23011 N23012 Segment
X23012 N23012 N23013 Segment
X23013 N23013 N23014 Segment
X23014 N23014 N23015 Segment
X23015 N23015 N23016 Segment
X23016 N23016 N23017 Segment
X23017 N23017 N23018 Segment
X23018 N23018 N23019 Segment
X23019 N23019 N23020 Segment
X23020 N23020 N23021 Segment
X23021 N23021 N23022 Segment
X23022 N23022 N23023 Segment
X23023 N23023 N23024 Segment
X23024 N23024 N23025 Segment
X23025 N23025 N23026 Segment
X23026 N23026 N23027 Segment
X23027 N23027 N23028 Segment
X23028 N23028 N23029 Segment
X23029 N23029 N23030 Segment
X23030 N23030 N23031 Segment
X23031 N23031 N23032 Segment
X23032 N23032 N23033 Segment
X23033 N23033 N23034 Segment
X23034 N23034 N23035 Segment
X23035 N23035 N23036 Segment
X23036 N23036 N23037 Segment
X23037 N23037 N23038 Segment
X23038 N23038 N23039 Segment
X23039 N23039 N23040 Segment
X23040 N23040 N23041 Segment
X23041 N23041 N23042 Segment
X23042 N23042 N23043 Segment
X23043 N23043 N23044 Segment
X23044 N23044 N23045 Segment
X23045 N23045 N23046 Segment
X23046 N23046 N23047 Segment
X23047 N23047 N23048 Segment
X23048 N23048 N23049 Segment
X23049 N23049 N23050 Segment
X23050 N23050 N23051 Segment
X23051 N23051 N23052 Segment
X23052 N23052 N23053 Segment
X23053 N23053 N23054 Segment
X23054 N23054 N23055 Segment
X23055 N23055 N23056 Segment
X23056 N23056 N23057 Segment
X23057 N23057 N23058 Segment
X23058 N23058 N23059 Segment
X23059 N23059 N23060 Segment
X23060 N23060 N23061 Segment
X23061 N23061 N23062 Segment
X23062 N23062 N23063 Segment
X23063 N23063 N23064 Segment
X23064 N23064 N23065 Segment
X23065 N23065 N23066 Segment
X23066 N23066 N23067 Segment
X23067 N23067 N23068 Segment
X23068 N23068 N23069 Segment
X23069 N23069 N23070 Segment
X23070 N23070 N23071 Segment
X23071 N23071 N23072 Segment
X23072 N23072 N23073 Segment
X23073 N23073 N23074 Segment
X23074 N23074 N23075 Segment
X23075 N23075 N23076 Segment
X23076 N23076 N23077 Segment
X23077 N23077 N23078 Segment
X23078 N23078 N23079 Segment
X23079 N23079 N23080 Segment
X23080 N23080 N23081 Segment
X23081 N23081 N23082 Segment
X23082 N23082 N23083 Segment
X23083 N23083 N23084 Segment
X23084 N23084 N23085 Segment
X23085 N23085 N23086 Segment
X23086 N23086 N23087 Segment
X23087 N23087 N23088 Segment
X23088 N23088 N23089 Segment
X23089 N23089 N23090 Segment
X23090 N23090 N23091 Segment
X23091 N23091 N23092 Segment
X23092 N23092 N23093 Segment
X23093 N23093 N23094 Segment
X23094 N23094 N23095 Segment
X23095 N23095 N23096 Segment
X23096 N23096 N23097 Segment
X23097 N23097 N23098 Segment
X23098 N23098 N23099 Segment
X23099 N23099 N23100 Segment
X23100 N23100 N23101 Segment
X23101 N23101 N23102 Segment
X23102 N23102 N23103 Segment
X23103 N23103 N23104 Segment
X23104 N23104 N23105 Segment
X23105 N23105 N23106 Segment
X23106 N23106 N23107 Segment
X23107 N23107 N23108 Segment
X23108 N23108 N23109 Segment
X23109 N23109 N23110 Segment
X23110 N23110 N23111 Segment
X23111 N23111 N23112 Segment
X23112 N23112 N23113 Segment
X23113 N23113 N23114 Segment
X23114 N23114 N23115 Segment
X23115 N23115 N23116 Segment
X23116 N23116 N23117 Segment
X23117 N23117 N23118 Segment
X23118 N23118 N23119 Segment
X23119 N23119 N23120 Segment
X23120 N23120 N23121 Segment
X23121 N23121 N23122 Segment
X23122 N23122 N23123 Segment
X23123 N23123 N23124 Segment
X23124 N23124 N23125 Segment
X23125 N23125 N23126 Segment
X23126 N23126 N23127 Segment
X23127 N23127 N23128 Segment
X23128 N23128 N23129 Segment
X23129 N23129 N23130 Segment
X23130 N23130 N23131 Segment
X23131 N23131 N23132 Segment
X23132 N23132 N23133 Segment
X23133 N23133 N23134 Segment
X23134 N23134 N23135 Segment
X23135 N23135 N23136 Segment
X23136 N23136 N23137 Segment
X23137 N23137 N23138 Segment
X23138 N23138 N23139 Segment
X23139 N23139 N23140 Segment
X23140 N23140 N23141 Segment
X23141 N23141 N23142 Segment
X23142 N23142 N23143 Segment
X23143 N23143 N23144 Segment
X23144 N23144 N23145 Segment
X23145 N23145 N23146 Segment
X23146 N23146 N23147 Segment
X23147 N23147 N23148 Segment
X23148 N23148 N23149 Segment
X23149 N23149 N23150 Segment
X23150 N23150 N23151 Segment
X23151 N23151 N23152 Segment
X23152 N23152 N23153 Segment
X23153 N23153 N23154 Segment
X23154 N23154 N23155 Segment
X23155 N23155 N23156 Segment
X23156 N23156 N23157 Segment
X23157 N23157 N23158 Segment
X23158 N23158 N23159 Segment
X23159 N23159 N23160 Segment
X23160 N23160 N23161 Segment
X23161 N23161 N23162 Segment
X23162 N23162 N23163 Segment
X23163 N23163 N23164 Segment
X23164 N23164 N23165 Segment
X23165 N23165 N23166 Segment
X23166 N23166 N23167 Segment
X23167 N23167 N23168 Segment
X23168 N23168 N23169 Segment
X23169 N23169 N23170 Segment
X23170 N23170 N23171 Segment
X23171 N23171 N23172 Segment
X23172 N23172 N23173 Segment
X23173 N23173 N23174 Segment
X23174 N23174 N23175 Segment
X23175 N23175 N23176 Segment
X23176 N23176 N23177 Segment
X23177 N23177 N23178 Segment
X23178 N23178 N23179 Segment
X23179 N23179 N23180 Segment
X23180 N23180 N23181 Segment
X23181 N23181 N23182 Segment
X23182 N23182 N23183 Segment
X23183 N23183 N23184 Segment
X23184 N23184 N23185 Segment
X23185 N23185 N23186 Segment
X23186 N23186 N23187 Segment
X23187 N23187 N23188 Segment
X23188 N23188 N23189 Segment
X23189 N23189 N23190 Segment
X23190 N23190 N23191 Segment
X23191 N23191 N23192 Segment
X23192 N23192 N23193 Segment
X23193 N23193 N23194 Segment
X23194 N23194 N23195 Segment
X23195 N23195 N23196 Segment
X23196 N23196 N23197 Segment
X23197 N23197 N23198 Segment
X23198 N23198 N23199 Segment
X23199 N23199 N23200 Segment
X23200 N23200 N23201 Segment
X23201 N23201 N23202 Segment
X23202 N23202 N23203 Segment
X23203 N23203 N23204 Segment
X23204 N23204 N23205 Segment
X23205 N23205 N23206 Segment
X23206 N23206 N23207 Segment
X23207 N23207 N23208 Segment
X23208 N23208 N23209 Segment
X23209 N23209 N23210 Segment
X23210 N23210 N23211 Segment
X23211 N23211 N23212 Segment
X23212 N23212 N23213 Segment
X23213 N23213 N23214 Segment
X23214 N23214 N23215 Segment
X23215 N23215 N23216 Segment
X23216 N23216 N23217 Segment
X23217 N23217 N23218 Segment
X23218 N23218 N23219 Segment
X23219 N23219 N23220 Segment
X23220 N23220 N23221 Segment
X23221 N23221 N23222 Segment
X23222 N23222 N23223 Segment
X23223 N23223 N23224 Segment
X23224 N23224 N23225 Segment
X23225 N23225 N23226 Segment
X23226 N23226 N23227 Segment
X23227 N23227 N23228 Segment
X23228 N23228 N23229 Segment
X23229 N23229 N23230 Segment
X23230 N23230 N23231 Segment
X23231 N23231 N23232 Segment
X23232 N23232 N23233 Segment
X23233 N23233 N23234 Segment
X23234 N23234 N23235 Segment
X23235 N23235 N23236 Segment
X23236 N23236 N23237 Segment
X23237 N23237 N23238 Segment
X23238 N23238 N23239 Segment
X23239 N23239 N23240 Segment
X23240 N23240 N23241 Segment
X23241 N23241 N23242 Segment
X23242 N23242 N23243 Segment
X23243 N23243 N23244 Segment
X23244 N23244 N23245 Segment
X23245 N23245 N23246 Segment
X23246 N23246 N23247 Segment
X23247 N23247 N23248 Segment
X23248 N23248 N23249 Segment
X23249 N23249 N23250 Segment
X23250 N23250 N23251 Segment
X23251 N23251 N23252 Segment
X23252 N23252 N23253 Segment
X23253 N23253 N23254 Segment
X23254 N23254 N23255 Segment
X23255 N23255 N23256 Segment
X23256 N23256 N23257 Segment
X23257 N23257 N23258 Segment
X23258 N23258 N23259 Segment
X23259 N23259 N23260 Segment
X23260 N23260 N23261 Segment
X23261 N23261 N23262 Segment
X23262 N23262 N23263 Segment
X23263 N23263 N23264 Segment
X23264 N23264 N23265 Segment
X23265 N23265 N23266 Segment
X23266 N23266 N23267 Segment
X23267 N23267 N23268 Segment
X23268 N23268 N23269 Segment
X23269 N23269 N23270 Segment
X23270 N23270 N23271 Segment
X23271 N23271 N23272 Segment
X23272 N23272 N23273 Segment
X23273 N23273 N23274 Segment
X23274 N23274 N23275 Segment
X23275 N23275 N23276 Segment
X23276 N23276 N23277 Segment
X23277 N23277 N23278 Segment
X23278 N23278 N23279 Segment
X23279 N23279 N23280 Segment
X23280 N23280 N23281 Segment
X23281 N23281 N23282 Segment
X23282 N23282 N23283 Segment
X23283 N23283 N23284 Segment
X23284 N23284 N23285 Segment
X23285 N23285 N23286 Segment
X23286 N23286 N23287 Segment
X23287 N23287 N23288 Segment
X23288 N23288 N23289 Segment
X23289 N23289 N23290 Segment
X23290 N23290 N23291 Segment
X23291 N23291 N23292 Segment
X23292 N23292 N23293 Segment
X23293 N23293 N23294 Segment
X23294 N23294 N23295 Segment
X23295 N23295 N23296 Segment
X23296 N23296 N23297 Segment
X23297 N23297 N23298 Segment
X23298 N23298 N23299 Segment
X23299 N23299 N23300 Segment
X23300 N23300 N23301 Segment
X23301 N23301 N23302 Segment
X23302 N23302 N23303 Segment
X23303 N23303 N23304 Segment
X23304 N23304 N23305 Segment
X23305 N23305 N23306 Segment
X23306 N23306 N23307 Segment
X23307 N23307 N23308 Segment
X23308 N23308 N23309 Segment
X23309 N23309 N23310 Segment
X23310 N23310 N23311 Segment
X23311 N23311 N23312 Segment
X23312 N23312 N23313 Segment
X23313 N23313 N23314 Segment
X23314 N23314 N23315 Segment
X23315 N23315 N23316 Segment
X23316 N23316 N23317 Segment
X23317 N23317 N23318 Segment
X23318 N23318 N23319 Segment
X23319 N23319 N23320 Segment
X23320 N23320 N23321 Segment
X23321 N23321 N23322 Segment
X23322 N23322 N23323 Segment
X23323 N23323 N23324 Segment
X23324 N23324 N23325 Segment
X23325 N23325 N23326 Segment
X23326 N23326 N23327 Segment
X23327 N23327 N23328 Segment
X23328 N23328 N23329 Segment
X23329 N23329 N23330 Segment
X23330 N23330 N23331 Segment
X23331 N23331 N23332 Segment
X23332 N23332 N23333 Segment
X23333 N23333 N23334 Segment
X23334 N23334 N23335 Segment
X23335 N23335 N23336 Segment
X23336 N23336 N23337 Segment
X23337 N23337 N23338 Segment
X23338 N23338 N23339 Segment
X23339 N23339 N23340 Segment
X23340 N23340 N23341 Segment
X23341 N23341 N23342 Segment
X23342 N23342 N23343 Segment
X23343 N23343 N23344 Segment
X23344 N23344 N23345 Segment
X23345 N23345 N23346 Segment
X23346 N23346 N23347 Segment
X23347 N23347 N23348 Segment
X23348 N23348 N23349 Segment
X23349 N23349 N23350 Segment
X23350 N23350 N23351 Segment
X23351 N23351 N23352 Segment
X23352 N23352 N23353 Segment
X23353 N23353 N23354 Segment
X23354 N23354 N23355 Segment
X23355 N23355 N23356 Segment
X23356 N23356 N23357 Segment
X23357 N23357 N23358 Segment
X23358 N23358 N23359 Segment
X23359 N23359 N23360 Segment
X23360 N23360 N23361 Segment
X23361 N23361 N23362 Segment
X23362 N23362 N23363 Segment
X23363 N23363 N23364 Segment
X23364 N23364 N23365 Segment
X23365 N23365 N23366 Segment
X23366 N23366 N23367 Segment
X23367 N23367 N23368 Segment
X23368 N23368 N23369 Segment
X23369 N23369 N23370 Segment
X23370 N23370 N23371 Segment
X23371 N23371 N23372 Segment
X23372 N23372 N23373 Segment
X23373 N23373 N23374 Segment
X23374 N23374 N23375 Segment
X23375 N23375 N23376 Segment
X23376 N23376 N23377 Segment
X23377 N23377 N23378 Segment
X23378 N23378 N23379 Segment
X23379 N23379 N23380 Segment
X23380 N23380 N23381 Segment
X23381 N23381 N23382 Segment
X23382 N23382 N23383 Segment
X23383 N23383 N23384 Segment
X23384 N23384 N23385 Segment
X23385 N23385 N23386 Segment
X23386 N23386 N23387 Segment
X23387 N23387 N23388 Segment
X23388 N23388 N23389 Segment
X23389 N23389 N23390 Segment
X23390 N23390 N23391 Segment
X23391 N23391 N23392 Segment
X23392 N23392 N23393 Segment
X23393 N23393 N23394 Segment
X23394 N23394 N23395 Segment
X23395 N23395 N23396 Segment
X23396 N23396 N23397 Segment
X23397 N23397 N23398 Segment
X23398 N23398 N23399 Segment
X23399 N23399 N23400 Segment
X23400 N23400 N23401 Segment
X23401 N23401 N23402 Segment
X23402 N23402 N23403 Segment
X23403 N23403 N23404 Segment
X23404 N23404 N23405 Segment
X23405 N23405 N23406 Segment
X23406 N23406 N23407 Segment
X23407 N23407 N23408 Segment
X23408 N23408 N23409 Segment
X23409 N23409 N23410 Segment
X23410 N23410 N23411 Segment
X23411 N23411 N23412 Segment
X23412 N23412 N23413 Segment
X23413 N23413 N23414 Segment
X23414 N23414 N23415 Segment
X23415 N23415 N23416 Segment
X23416 N23416 N23417 Segment
X23417 N23417 N23418 Segment
X23418 N23418 N23419 Segment
X23419 N23419 N23420 Segment
X23420 N23420 N23421 Segment
X23421 N23421 N23422 Segment
X23422 N23422 N23423 Segment
X23423 N23423 N23424 Segment
X23424 N23424 N23425 Segment
X23425 N23425 N23426 Segment
X23426 N23426 N23427 Segment
X23427 N23427 N23428 Segment
X23428 N23428 N23429 Segment
X23429 N23429 N23430 Segment
X23430 N23430 N23431 Segment
X23431 N23431 N23432 Segment
X23432 N23432 N23433 Segment
X23433 N23433 N23434 Segment
X23434 N23434 N23435 Segment
X23435 N23435 N23436 Segment
X23436 N23436 N23437 Segment
X23437 N23437 N23438 Segment
X23438 N23438 N23439 Segment
X23439 N23439 N23440 Segment
X23440 N23440 N23441 Segment
X23441 N23441 N23442 Segment
X23442 N23442 N23443 Segment
X23443 N23443 N23444 Segment
X23444 N23444 N23445 Segment
X23445 N23445 N23446 Segment
X23446 N23446 N23447 Segment
X23447 N23447 N23448 Segment
X23448 N23448 N23449 Segment
X23449 N23449 N23450 Segment
X23450 N23450 N23451 Segment
X23451 N23451 N23452 Segment
X23452 N23452 N23453 Segment
X23453 N23453 N23454 Segment
X23454 N23454 N23455 Segment
X23455 N23455 N23456 Segment
X23456 N23456 N23457 Segment
X23457 N23457 N23458 Segment
X23458 N23458 N23459 Segment
X23459 N23459 N23460 Segment
X23460 N23460 N23461 Segment
X23461 N23461 N23462 Segment
X23462 N23462 N23463 Segment
X23463 N23463 N23464 Segment
X23464 N23464 N23465 Segment
X23465 N23465 N23466 Segment
X23466 N23466 N23467 Segment
X23467 N23467 N23468 Segment
X23468 N23468 N23469 Segment
X23469 N23469 N23470 Segment
X23470 N23470 N23471 Segment
X23471 N23471 N23472 Segment
X23472 N23472 N23473 Segment
X23473 N23473 N23474 Segment
X23474 N23474 N23475 Segment
X23475 N23475 N23476 Segment
X23476 N23476 N23477 Segment
X23477 N23477 N23478 Segment
X23478 N23478 N23479 Segment
X23479 N23479 N23480 Segment
X23480 N23480 N23481 Segment
X23481 N23481 N23482 Segment
X23482 N23482 N23483 Segment
X23483 N23483 N23484 Segment
X23484 N23484 N23485 Segment
X23485 N23485 N23486 Segment
X23486 N23486 N23487 Segment
X23487 N23487 N23488 Segment
X23488 N23488 N23489 Segment
X23489 N23489 N23490 Segment
X23490 N23490 N23491 Segment
X23491 N23491 N23492 Segment
X23492 N23492 N23493 Segment
X23493 N23493 N23494 Segment
X23494 N23494 N23495 Segment
X23495 N23495 N23496 Segment
X23496 N23496 N23497 Segment
X23497 N23497 N23498 Segment
X23498 N23498 N23499 Segment
X23499 N23499 N23500 Segment
X23500 N23500 N23501 Segment
X23501 N23501 N23502 Segment
X23502 N23502 N23503 Segment
X23503 N23503 N23504 Segment
X23504 N23504 N23505 Segment
X23505 N23505 N23506 Segment
X23506 N23506 N23507 Segment
X23507 N23507 N23508 Segment
X23508 N23508 N23509 Segment
X23509 N23509 N23510 Segment
X23510 N23510 N23511 Segment
X23511 N23511 N23512 Segment
X23512 N23512 N23513 Segment
X23513 N23513 N23514 Segment
X23514 N23514 N23515 Segment
X23515 N23515 N23516 Segment
X23516 N23516 N23517 Segment
X23517 N23517 N23518 Segment
X23518 N23518 N23519 Segment
X23519 N23519 N23520 Segment
X23520 N23520 N23521 Segment
X23521 N23521 N23522 Segment
X23522 N23522 N23523 Segment
X23523 N23523 N23524 Segment
X23524 N23524 N23525 Segment
X23525 N23525 N23526 Segment
X23526 N23526 N23527 Segment
X23527 N23527 N23528 Segment
X23528 N23528 N23529 Segment
X23529 N23529 N23530 Segment
X23530 N23530 N23531 Segment
X23531 N23531 N23532 Segment
X23532 N23532 N23533 Segment
X23533 N23533 N23534 Segment
X23534 N23534 N23535 Segment
X23535 N23535 N23536 Segment
X23536 N23536 N23537 Segment
X23537 N23537 N23538 Segment
X23538 N23538 N23539 Segment
X23539 N23539 N23540 Segment
X23540 N23540 N23541 Segment
X23541 N23541 N23542 Segment
X23542 N23542 N23543 Segment
X23543 N23543 N23544 Segment
X23544 N23544 N23545 Segment
X23545 N23545 N23546 Segment
X23546 N23546 N23547 Segment
X23547 N23547 N23548 Segment
X23548 N23548 N23549 Segment
X23549 N23549 N23550 Segment
X23550 N23550 N23551 Segment
X23551 N23551 N23552 Segment
X23552 N23552 N23553 Segment
X23553 N23553 N23554 Segment
X23554 N23554 N23555 Segment
X23555 N23555 N23556 Segment
X23556 N23556 N23557 Segment
X23557 N23557 N23558 Segment
X23558 N23558 N23559 Segment
X23559 N23559 N23560 Segment
X23560 N23560 N23561 Segment
X23561 N23561 N23562 Segment
X23562 N23562 N23563 Segment
X23563 N23563 N23564 Segment
X23564 N23564 N23565 Segment
X23565 N23565 N23566 Segment
X23566 N23566 N23567 Segment
X23567 N23567 N23568 Segment
X23568 N23568 N23569 Segment
X23569 N23569 N23570 Segment
X23570 N23570 N23571 Segment
X23571 N23571 N23572 Segment
X23572 N23572 N23573 Segment
X23573 N23573 N23574 Segment
X23574 N23574 N23575 Segment
X23575 N23575 N23576 Segment
X23576 N23576 N23577 Segment
X23577 N23577 N23578 Segment
X23578 N23578 N23579 Segment
X23579 N23579 N23580 Segment
X23580 N23580 N23581 Segment
X23581 N23581 N23582 Segment
X23582 N23582 N23583 Segment
X23583 N23583 N23584 Segment
X23584 N23584 N23585 Segment
X23585 N23585 N23586 Segment
X23586 N23586 N23587 Segment
X23587 N23587 N23588 Segment
X23588 N23588 N23589 Segment
X23589 N23589 N23590 Segment
X23590 N23590 N23591 Segment
X23591 N23591 N23592 Segment
X23592 N23592 N23593 Segment
X23593 N23593 N23594 Segment
X23594 N23594 N23595 Segment
X23595 N23595 N23596 Segment
X23596 N23596 N23597 Segment
X23597 N23597 N23598 Segment
X23598 N23598 N23599 Segment
X23599 N23599 N23600 Segment
X23600 N23600 N23601 Segment
X23601 N23601 N23602 Segment
X23602 N23602 N23603 Segment
X23603 N23603 N23604 Segment
X23604 N23604 N23605 Segment
X23605 N23605 N23606 Segment
X23606 N23606 N23607 Segment
X23607 N23607 N23608 Segment
X23608 N23608 N23609 Segment
X23609 N23609 N23610 Segment
X23610 N23610 N23611 Segment
X23611 N23611 N23612 Segment
X23612 N23612 N23613 Segment
X23613 N23613 N23614 Segment
X23614 N23614 N23615 Segment
X23615 N23615 N23616 Segment
X23616 N23616 N23617 Segment
X23617 N23617 N23618 Segment
X23618 N23618 N23619 Segment
X23619 N23619 N23620 Segment
X23620 N23620 N23621 Segment
X23621 N23621 N23622 Segment
X23622 N23622 N23623 Segment
X23623 N23623 N23624 Segment
X23624 N23624 N23625 Segment
X23625 N23625 N23626 Segment
X23626 N23626 N23627 Segment
X23627 N23627 N23628 Segment
X23628 N23628 N23629 Segment
X23629 N23629 N23630 Segment
X23630 N23630 N23631 Segment
X23631 N23631 N23632 Segment
X23632 N23632 N23633 Segment
X23633 N23633 N23634 Segment
X23634 N23634 N23635 Segment
X23635 N23635 N23636 Segment
X23636 N23636 N23637 Segment
X23637 N23637 N23638 Segment
X23638 N23638 N23639 Segment
X23639 N23639 N23640 Segment
X23640 N23640 N23641 Segment
X23641 N23641 N23642 Segment
X23642 N23642 N23643 Segment
X23643 N23643 N23644 Segment
X23644 N23644 N23645 Segment
X23645 N23645 N23646 Segment
X23646 N23646 N23647 Segment
X23647 N23647 N23648 Segment
X23648 N23648 N23649 Segment
X23649 N23649 N23650 Segment
X23650 N23650 N23651 Segment
X23651 N23651 N23652 Segment
X23652 N23652 N23653 Segment
X23653 N23653 N23654 Segment
X23654 N23654 N23655 Segment
X23655 N23655 N23656 Segment
X23656 N23656 N23657 Segment
X23657 N23657 N23658 Segment
X23658 N23658 N23659 Segment
X23659 N23659 N23660 Segment
X23660 N23660 N23661 Segment
X23661 N23661 N23662 Segment
X23662 N23662 N23663 Segment
X23663 N23663 N23664 Segment
X23664 N23664 N23665 Segment
X23665 N23665 N23666 Segment
X23666 N23666 N23667 Segment
X23667 N23667 N23668 Segment
X23668 N23668 N23669 Segment
X23669 N23669 N23670 Segment
X23670 N23670 N23671 Segment
X23671 N23671 N23672 Segment
X23672 N23672 N23673 Segment
X23673 N23673 N23674 Segment
X23674 N23674 N23675 Segment
X23675 N23675 N23676 Segment
X23676 N23676 N23677 Segment
X23677 N23677 N23678 Segment
X23678 N23678 N23679 Segment
X23679 N23679 N23680 Segment
X23680 N23680 N23681 Segment
X23681 N23681 N23682 Segment
X23682 N23682 N23683 Segment
X23683 N23683 N23684 Segment
X23684 N23684 N23685 Segment
X23685 N23685 N23686 Segment
X23686 N23686 N23687 Segment
X23687 N23687 N23688 Segment
X23688 N23688 N23689 Segment
X23689 N23689 N23690 Segment
X23690 N23690 N23691 Segment
X23691 N23691 N23692 Segment
X23692 N23692 N23693 Segment
X23693 N23693 N23694 Segment
X23694 N23694 N23695 Segment
X23695 N23695 N23696 Segment
X23696 N23696 N23697 Segment
X23697 N23697 N23698 Segment
X23698 N23698 N23699 Segment
X23699 N23699 N23700 Segment
X23700 N23700 N23701 Segment
X23701 N23701 N23702 Segment
X23702 N23702 N23703 Segment
X23703 N23703 N23704 Segment
X23704 N23704 N23705 Segment
X23705 N23705 N23706 Segment
X23706 N23706 N23707 Segment
X23707 N23707 N23708 Segment
X23708 N23708 N23709 Segment
X23709 N23709 N23710 Segment
X23710 N23710 N23711 Segment
X23711 N23711 N23712 Segment
X23712 N23712 N23713 Segment
X23713 N23713 N23714 Segment
X23714 N23714 N23715 Segment
X23715 N23715 N23716 Segment
X23716 N23716 N23717 Segment
X23717 N23717 N23718 Segment
X23718 N23718 N23719 Segment
X23719 N23719 N23720 Segment
X23720 N23720 N23721 Segment
X23721 N23721 N23722 Segment
X23722 N23722 N23723 Segment
X23723 N23723 N23724 Segment
X23724 N23724 N23725 Segment
X23725 N23725 N23726 Segment
X23726 N23726 N23727 Segment
X23727 N23727 N23728 Segment
X23728 N23728 N23729 Segment
X23729 N23729 N23730 Segment
X23730 N23730 N23731 Segment
X23731 N23731 N23732 Segment
X23732 N23732 N23733 Segment
X23733 N23733 N23734 Segment
X23734 N23734 N23735 Segment
X23735 N23735 N23736 Segment
X23736 N23736 N23737 Segment
X23737 N23737 N23738 Segment
X23738 N23738 N23739 Segment
X23739 N23739 N23740 Segment
X23740 N23740 N23741 Segment
X23741 N23741 N23742 Segment
X23742 N23742 N23743 Segment
X23743 N23743 N23744 Segment
X23744 N23744 N23745 Segment
X23745 N23745 N23746 Segment
X23746 N23746 N23747 Segment
X23747 N23747 N23748 Segment
X23748 N23748 N23749 Segment
X23749 N23749 N23750 Segment
X23750 N23750 N23751 Segment
X23751 N23751 N23752 Segment
X23752 N23752 N23753 Segment
X23753 N23753 N23754 Segment
X23754 N23754 N23755 Segment
X23755 N23755 N23756 Segment
X23756 N23756 N23757 Segment
X23757 N23757 N23758 Segment
X23758 N23758 N23759 Segment
X23759 N23759 N23760 Segment
X23760 N23760 N23761 Segment
X23761 N23761 N23762 Segment
X23762 N23762 N23763 Segment
X23763 N23763 N23764 Segment
X23764 N23764 N23765 Segment
X23765 N23765 N23766 Segment
X23766 N23766 N23767 Segment
X23767 N23767 N23768 Segment
X23768 N23768 N23769 Segment
X23769 N23769 N23770 Segment
X23770 N23770 N23771 Segment
X23771 N23771 N23772 Segment
X23772 N23772 N23773 Segment
X23773 N23773 N23774 Segment
X23774 N23774 N23775 Segment
X23775 N23775 N23776 Segment
X23776 N23776 N23777 Segment
X23777 N23777 N23778 Segment
X23778 N23778 N23779 Segment
X23779 N23779 N23780 Segment
X23780 N23780 N23781 Segment
X23781 N23781 N23782 Segment
X23782 N23782 N23783 Segment
X23783 N23783 N23784 Segment
X23784 N23784 N23785 Segment
X23785 N23785 N23786 Segment
X23786 N23786 N23787 Segment
X23787 N23787 N23788 Segment
X23788 N23788 N23789 Segment
X23789 N23789 N23790 Segment
X23790 N23790 N23791 Segment
X23791 N23791 N23792 Segment
X23792 N23792 N23793 Segment
X23793 N23793 N23794 Segment
X23794 N23794 N23795 Segment
X23795 N23795 N23796 Segment
X23796 N23796 N23797 Segment
X23797 N23797 N23798 Segment
X23798 N23798 N23799 Segment
X23799 N23799 N23800 Segment
X23800 N23800 N23801 Segment
X23801 N23801 N23802 Segment
X23802 N23802 N23803 Segment
X23803 N23803 N23804 Segment
X23804 N23804 N23805 Segment
X23805 N23805 N23806 Segment
X23806 N23806 N23807 Segment
X23807 N23807 N23808 Segment
X23808 N23808 N23809 Segment
X23809 N23809 N23810 Segment
X23810 N23810 N23811 Segment
X23811 N23811 N23812 Segment
X23812 N23812 N23813 Segment
X23813 N23813 N23814 Segment
X23814 N23814 N23815 Segment
X23815 N23815 N23816 Segment
X23816 N23816 N23817 Segment
X23817 N23817 N23818 Segment
X23818 N23818 N23819 Segment
X23819 N23819 N23820 Segment
X23820 N23820 N23821 Segment
X23821 N23821 N23822 Segment
X23822 N23822 N23823 Segment
X23823 N23823 N23824 Segment
X23824 N23824 N23825 Segment
X23825 N23825 N23826 Segment
X23826 N23826 N23827 Segment
X23827 N23827 N23828 Segment
X23828 N23828 N23829 Segment
X23829 N23829 N23830 Segment
X23830 N23830 N23831 Segment
X23831 N23831 N23832 Segment
X23832 N23832 N23833 Segment
X23833 N23833 N23834 Segment
X23834 N23834 N23835 Segment
X23835 N23835 N23836 Segment
X23836 N23836 N23837 Segment
X23837 N23837 N23838 Segment
X23838 N23838 N23839 Segment
X23839 N23839 N23840 Segment
X23840 N23840 N23841 Segment
X23841 N23841 N23842 Segment
X23842 N23842 N23843 Segment
X23843 N23843 N23844 Segment
X23844 N23844 N23845 Segment
X23845 N23845 N23846 Segment
X23846 N23846 N23847 Segment
X23847 N23847 N23848 Segment
X23848 N23848 N23849 Segment
X23849 N23849 N23850 Segment
X23850 N23850 N23851 Segment
X23851 N23851 N23852 Segment
X23852 N23852 N23853 Segment
X23853 N23853 N23854 Segment
X23854 N23854 N23855 Segment
X23855 N23855 N23856 Segment
X23856 N23856 N23857 Segment
X23857 N23857 N23858 Segment
X23858 N23858 N23859 Segment
X23859 N23859 N23860 Segment
X23860 N23860 N23861 Segment
X23861 N23861 N23862 Segment
X23862 N23862 N23863 Segment
X23863 N23863 N23864 Segment
X23864 N23864 N23865 Segment
X23865 N23865 N23866 Segment
X23866 N23866 N23867 Segment
X23867 N23867 N23868 Segment
X23868 N23868 N23869 Segment
X23869 N23869 N23870 Segment
X23870 N23870 N23871 Segment
X23871 N23871 N23872 Segment
X23872 N23872 N23873 Segment
X23873 N23873 N23874 Segment
X23874 N23874 N23875 Segment
X23875 N23875 N23876 Segment
X23876 N23876 N23877 Segment
X23877 N23877 N23878 Segment
X23878 N23878 N23879 Segment
X23879 N23879 N23880 Segment
X23880 N23880 N23881 Segment
X23881 N23881 N23882 Segment
X23882 N23882 N23883 Segment
X23883 N23883 N23884 Segment
X23884 N23884 N23885 Segment
X23885 N23885 N23886 Segment
X23886 N23886 N23887 Segment
X23887 N23887 N23888 Segment
X23888 N23888 N23889 Segment
X23889 N23889 N23890 Segment
X23890 N23890 N23891 Segment
X23891 N23891 N23892 Segment
X23892 N23892 N23893 Segment
X23893 N23893 N23894 Segment
X23894 N23894 N23895 Segment
X23895 N23895 N23896 Segment
X23896 N23896 N23897 Segment
X23897 N23897 N23898 Segment
X23898 N23898 N23899 Segment
X23899 N23899 N23900 Segment
X23900 N23900 N23901 Segment
X23901 N23901 N23902 Segment
X23902 N23902 N23903 Segment
X23903 N23903 N23904 Segment
X23904 N23904 N23905 Segment
X23905 N23905 N23906 Segment
X23906 N23906 N23907 Segment
X23907 N23907 N23908 Segment
X23908 N23908 N23909 Segment
X23909 N23909 N23910 Segment
X23910 N23910 N23911 Segment
X23911 N23911 N23912 Segment
X23912 N23912 N23913 Segment
X23913 N23913 N23914 Segment
X23914 N23914 N23915 Segment
X23915 N23915 N23916 Segment
X23916 N23916 N23917 Segment
X23917 N23917 N23918 Segment
X23918 N23918 N23919 Segment
X23919 N23919 N23920 Segment
X23920 N23920 N23921 Segment
X23921 N23921 N23922 Segment
X23922 N23922 N23923 Segment
X23923 N23923 N23924 Segment
X23924 N23924 N23925 Segment
X23925 N23925 N23926 Segment
X23926 N23926 N23927 Segment
X23927 N23927 N23928 Segment
X23928 N23928 N23929 Segment
X23929 N23929 N23930 Segment
X23930 N23930 N23931 Segment
X23931 N23931 N23932 Segment
X23932 N23932 N23933 Segment
X23933 N23933 N23934 Segment
X23934 N23934 N23935 Segment
X23935 N23935 N23936 Segment
X23936 N23936 N23937 Segment
X23937 N23937 N23938 Segment
X23938 N23938 N23939 Segment
X23939 N23939 N23940 Segment
X23940 N23940 N23941 Segment
X23941 N23941 N23942 Segment
X23942 N23942 N23943 Segment
X23943 N23943 N23944 Segment
X23944 N23944 N23945 Segment
X23945 N23945 N23946 Segment
X23946 N23946 N23947 Segment
X23947 N23947 N23948 Segment
X23948 N23948 N23949 Segment
X23949 N23949 N23950 Segment
X23950 N23950 N23951 Segment
X23951 N23951 N23952 Segment
X23952 N23952 N23953 Segment
X23953 N23953 N23954 Segment
X23954 N23954 N23955 Segment
X23955 N23955 N23956 Segment
X23956 N23956 N23957 Segment
X23957 N23957 N23958 Segment
X23958 N23958 N23959 Segment
X23959 N23959 N23960 Segment
X23960 N23960 N23961 Segment
X23961 N23961 N23962 Segment
X23962 N23962 N23963 Segment
X23963 N23963 N23964 Segment
X23964 N23964 N23965 Segment
X23965 N23965 N23966 Segment
X23966 N23966 N23967 Segment
X23967 N23967 N23968 Segment
X23968 N23968 N23969 Segment
X23969 N23969 N23970 Segment
X23970 N23970 N23971 Segment
X23971 N23971 N23972 Segment
X23972 N23972 N23973 Segment
X23973 N23973 N23974 Segment
X23974 N23974 N23975 Segment
X23975 N23975 N23976 Segment
X23976 N23976 N23977 Segment
X23977 N23977 N23978 Segment
X23978 N23978 N23979 Segment
X23979 N23979 N23980 Segment
X23980 N23980 N23981 Segment
X23981 N23981 N23982 Segment
X23982 N23982 N23983 Segment
X23983 N23983 N23984 Segment
X23984 N23984 N23985 Segment
X23985 N23985 N23986 Segment
X23986 N23986 N23987 Segment
X23987 N23987 N23988 Segment
X23988 N23988 N23989 Segment
X23989 N23989 N23990 Segment
X23990 N23990 N23991 Segment
X23991 N23991 N23992 Segment
X23992 N23992 N23993 Segment
X23993 N23993 N23994 Segment
X23994 N23994 N23995 Segment
X23995 N23995 N23996 Segment
X23996 N23996 N23997 Segment
X23997 N23997 N23998 Segment
X23998 N23998 N23999 Segment
X23999 N23999 N24000 Segment
X24000 N24000 N24001 Segment
X24001 N24001 N24002 Segment
X24002 N24002 N24003 Segment
X24003 N24003 N24004 Segment
X24004 N24004 N24005 Segment
X24005 N24005 N24006 Segment
X24006 N24006 N24007 Segment
X24007 N24007 N24008 Segment
X24008 N24008 N24009 Segment
X24009 N24009 N24010 Segment
X24010 N24010 N24011 Segment
X24011 N24011 N24012 Segment
X24012 N24012 N24013 Segment
X24013 N24013 N24014 Segment
X24014 N24014 N24015 Segment
X24015 N24015 N24016 Segment
X24016 N24016 N24017 Segment
X24017 N24017 N24018 Segment
X24018 N24018 N24019 Segment
X24019 N24019 N24020 Segment
X24020 N24020 N24021 Segment
X24021 N24021 N24022 Segment
X24022 N24022 N24023 Segment
X24023 N24023 N24024 Segment
X24024 N24024 N24025 Segment
X24025 N24025 N24026 Segment
X24026 N24026 N24027 Segment
X24027 N24027 N24028 Segment
X24028 N24028 N24029 Segment
X24029 N24029 N24030 Segment
X24030 N24030 N24031 Segment
X24031 N24031 N24032 Segment
X24032 N24032 N24033 Segment
X24033 N24033 N24034 Segment
X24034 N24034 N24035 Segment
X24035 N24035 N24036 Segment
X24036 N24036 N24037 Segment
X24037 N24037 N24038 Segment
X24038 N24038 N24039 Segment
X24039 N24039 N24040 Segment
X24040 N24040 N24041 Segment
X24041 N24041 N24042 Segment
X24042 N24042 N24043 Segment
X24043 N24043 N24044 Segment
X24044 N24044 N24045 Segment
X24045 N24045 N24046 Segment
X24046 N24046 N24047 Segment
X24047 N24047 N24048 Segment
X24048 N24048 N24049 Segment
X24049 N24049 N24050 Segment
X24050 N24050 N24051 Segment
X24051 N24051 N24052 Segment
X24052 N24052 N24053 Segment
X24053 N24053 N24054 Segment
X24054 N24054 N24055 Segment
X24055 N24055 N24056 Segment
X24056 N24056 N24057 Segment
X24057 N24057 N24058 Segment
X24058 N24058 N24059 Segment
X24059 N24059 N24060 Segment
X24060 N24060 N24061 Segment
X24061 N24061 N24062 Segment
X24062 N24062 N24063 Segment
X24063 N24063 N24064 Segment
X24064 N24064 N24065 Segment
X24065 N24065 N24066 Segment
X24066 N24066 N24067 Segment
X24067 N24067 N24068 Segment
X24068 N24068 N24069 Segment
X24069 N24069 N24070 Segment
X24070 N24070 N24071 Segment
X24071 N24071 N24072 Segment
X24072 N24072 N24073 Segment
X24073 N24073 N24074 Segment
X24074 N24074 N24075 Segment
X24075 N24075 N24076 Segment
X24076 N24076 N24077 Segment
X24077 N24077 N24078 Segment
X24078 N24078 N24079 Segment
X24079 N24079 N24080 Segment
X24080 N24080 N24081 Segment
X24081 N24081 N24082 Segment
X24082 N24082 N24083 Segment
X24083 N24083 N24084 Segment
X24084 N24084 N24085 Segment
X24085 N24085 N24086 Segment
X24086 N24086 N24087 Segment
X24087 N24087 N24088 Segment
X24088 N24088 N24089 Segment
X24089 N24089 N24090 Segment
X24090 N24090 N24091 Segment
X24091 N24091 N24092 Segment
X24092 N24092 N24093 Segment
X24093 N24093 N24094 Segment
X24094 N24094 N24095 Segment
X24095 N24095 N24096 Segment
X24096 N24096 N24097 Segment
X24097 N24097 N24098 Segment
X24098 N24098 N24099 Segment
X24099 N24099 N24100 Segment
X24100 N24100 N24101 Segment
X24101 N24101 N24102 Segment
X24102 N24102 N24103 Segment
X24103 N24103 N24104 Segment
X24104 N24104 N24105 Segment
X24105 N24105 N24106 Segment
X24106 N24106 N24107 Segment
X24107 N24107 N24108 Segment
X24108 N24108 N24109 Segment
X24109 N24109 N24110 Segment
X24110 N24110 N24111 Segment
X24111 N24111 N24112 Segment
X24112 N24112 N24113 Segment
X24113 N24113 N24114 Segment
X24114 N24114 N24115 Segment
X24115 N24115 N24116 Segment
X24116 N24116 N24117 Segment
X24117 N24117 N24118 Segment
X24118 N24118 N24119 Segment
X24119 N24119 N24120 Segment
X24120 N24120 N24121 Segment
X24121 N24121 N24122 Segment
X24122 N24122 N24123 Segment
X24123 N24123 N24124 Segment
X24124 N24124 N24125 Segment
X24125 N24125 N24126 Segment
X24126 N24126 N24127 Segment
X24127 N24127 N24128 Segment
X24128 N24128 N24129 Segment
X24129 N24129 N24130 Segment
X24130 N24130 N24131 Segment
X24131 N24131 N24132 Segment
X24132 N24132 N24133 Segment
X24133 N24133 N24134 Segment
X24134 N24134 N24135 Segment
X24135 N24135 N24136 Segment
X24136 N24136 N24137 Segment
X24137 N24137 N24138 Segment
X24138 N24138 N24139 Segment
X24139 N24139 N24140 Segment
X24140 N24140 N24141 Segment
X24141 N24141 N24142 Segment
X24142 N24142 N24143 Segment
X24143 N24143 N24144 Segment
X24144 N24144 N24145 Segment
X24145 N24145 N24146 Segment
X24146 N24146 N24147 Segment
X24147 N24147 N24148 Segment
X24148 N24148 N24149 Segment
X24149 N24149 N24150 Segment
X24150 N24150 N24151 Segment
X24151 N24151 N24152 Segment
X24152 N24152 N24153 Segment
X24153 N24153 N24154 Segment
X24154 N24154 N24155 Segment
X24155 N24155 N24156 Segment
X24156 N24156 N24157 Segment
X24157 N24157 N24158 Segment
X24158 N24158 N24159 Segment
X24159 N24159 N24160 Segment
X24160 N24160 N24161 Segment
X24161 N24161 N24162 Segment
X24162 N24162 N24163 Segment
X24163 N24163 N24164 Segment
X24164 N24164 N24165 Segment
X24165 N24165 N24166 Segment
X24166 N24166 N24167 Segment
X24167 N24167 N24168 Segment
X24168 N24168 N24169 Segment
X24169 N24169 N24170 Segment
X24170 N24170 N24171 Segment
X24171 N24171 N24172 Segment
X24172 N24172 N24173 Segment
X24173 N24173 N24174 Segment
X24174 N24174 N24175 Segment
X24175 N24175 N24176 Segment
X24176 N24176 N24177 Segment
X24177 N24177 N24178 Segment
X24178 N24178 N24179 Segment
X24179 N24179 N24180 Segment
X24180 N24180 N24181 Segment
X24181 N24181 N24182 Segment
X24182 N24182 N24183 Segment
X24183 N24183 N24184 Segment
X24184 N24184 N24185 Segment
X24185 N24185 N24186 Segment
X24186 N24186 N24187 Segment
X24187 N24187 N24188 Segment
X24188 N24188 N24189 Segment
X24189 N24189 N24190 Segment
X24190 N24190 N24191 Segment
X24191 N24191 N24192 Segment
X24192 N24192 N24193 Segment
X24193 N24193 N24194 Segment
X24194 N24194 N24195 Segment
X24195 N24195 N24196 Segment
X24196 N24196 N24197 Segment
X24197 N24197 N24198 Segment
X24198 N24198 N24199 Segment
X24199 N24199 N24200 Segment
X24200 N24200 N24201 Segment
X24201 N24201 N24202 Segment
X24202 N24202 N24203 Segment
X24203 N24203 N24204 Segment
X24204 N24204 N24205 Segment
X24205 N24205 N24206 Segment
X24206 N24206 N24207 Segment
X24207 N24207 N24208 Segment
X24208 N24208 N24209 Segment
X24209 N24209 N24210 Segment
X24210 N24210 N24211 Segment
X24211 N24211 N24212 Segment
X24212 N24212 N24213 Segment
X24213 N24213 N24214 Segment
X24214 N24214 N24215 Segment
X24215 N24215 N24216 Segment
X24216 N24216 N24217 Segment
X24217 N24217 N24218 Segment
X24218 N24218 N24219 Segment
X24219 N24219 N24220 Segment
X24220 N24220 N24221 Segment
X24221 N24221 N24222 Segment
X24222 N24222 N24223 Segment
X24223 N24223 N24224 Segment
X24224 N24224 N24225 Segment
X24225 N24225 N24226 Segment
X24226 N24226 N24227 Segment
X24227 N24227 N24228 Segment
X24228 N24228 N24229 Segment
X24229 N24229 N24230 Segment
X24230 N24230 N24231 Segment
X24231 N24231 N24232 Segment
X24232 N24232 N24233 Segment
X24233 N24233 N24234 Segment
X24234 N24234 N24235 Segment
X24235 N24235 N24236 Segment
X24236 N24236 N24237 Segment
X24237 N24237 N24238 Segment
X24238 N24238 N24239 Segment
X24239 N24239 N24240 Segment
X24240 N24240 N24241 Segment
X24241 N24241 N24242 Segment
X24242 N24242 N24243 Segment
X24243 N24243 N24244 Segment
X24244 N24244 N24245 Segment
X24245 N24245 N24246 Segment
X24246 N24246 N24247 Segment
X24247 N24247 N24248 Segment
X24248 N24248 N24249 Segment
X24249 N24249 N24250 Segment
X24250 N24250 N24251 Segment
X24251 N24251 N24252 Segment
X24252 N24252 N24253 Segment
X24253 N24253 N24254 Segment
X24254 N24254 N24255 Segment
X24255 N24255 N24256 Segment
X24256 N24256 N24257 Segment
X24257 N24257 N24258 Segment
X24258 N24258 N24259 Segment
X24259 N24259 N24260 Segment
X24260 N24260 N24261 Segment
X24261 N24261 N24262 Segment
X24262 N24262 N24263 Segment
X24263 N24263 N24264 Segment
X24264 N24264 N24265 Segment
X24265 N24265 N24266 Segment
X24266 N24266 N24267 Segment
X24267 N24267 N24268 Segment
X24268 N24268 N24269 Segment
X24269 N24269 N24270 Segment
X24270 N24270 N24271 Segment
X24271 N24271 N24272 Segment
X24272 N24272 N24273 Segment
X24273 N24273 N24274 Segment
X24274 N24274 N24275 Segment
X24275 N24275 N24276 Segment
X24276 N24276 N24277 Segment
X24277 N24277 N24278 Segment
X24278 N24278 N24279 Segment
X24279 N24279 N24280 Segment
X24280 N24280 N24281 Segment
X24281 N24281 N24282 Segment
X24282 N24282 N24283 Segment
X24283 N24283 N24284 Segment
X24284 N24284 N24285 Segment
X24285 N24285 N24286 Segment
X24286 N24286 N24287 Segment
X24287 N24287 N24288 Segment
X24288 N24288 N24289 Segment
X24289 N24289 N24290 Segment
X24290 N24290 N24291 Segment
X24291 N24291 N24292 Segment
X24292 N24292 N24293 Segment
X24293 N24293 N24294 Segment
X24294 N24294 N24295 Segment
X24295 N24295 N24296 Segment
X24296 N24296 N24297 Segment
X24297 N24297 N24298 Segment
X24298 N24298 N24299 Segment
X24299 N24299 N24300 Segment
X24300 N24300 N24301 Segment
X24301 N24301 N24302 Segment
X24302 N24302 N24303 Segment
X24303 N24303 N24304 Segment
X24304 N24304 N24305 Segment
X24305 N24305 N24306 Segment
X24306 N24306 N24307 Segment
X24307 N24307 N24308 Segment
X24308 N24308 N24309 Segment
X24309 N24309 N24310 Segment
X24310 N24310 N24311 Segment
X24311 N24311 N24312 Segment
X24312 N24312 N24313 Segment
X24313 N24313 N24314 Segment
X24314 N24314 N24315 Segment
X24315 N24315 N24316 Segment
X24316 N24316 N24317 Segment
X24317 N24317 N24318 Segment
X24318 N24318 N24319 Segment
X24319 N24319 N24320 Segment
X24320 N24320 N24321 Segment
X24321 N24321 N24322 Segment
X24322 N24322 N24323 Segment
X24323 N24323 N24324 Segment
X24324 N24324 N24325 Segment
X24325 N24325 N24326 Segment
X24326 N24326 N24327 Segment
X24327 N24327 N24328 Segment
X24328 N24328 N24329 Segment
X24329 N24329 N24330 Segment
X24330 N24330 N24331 Segment
X24331 N24331 N24332 Segment
X24332 N24332 N24333 Segment
X24333 N24333 N24334 Segment
X24334 N24334 N24335 Segment
X24335 N24335 N24336 Segment
X24336 N24336 N24337 Segment
X24337 N24337 N24338 Segment
X24338 N24338 N24339 Segment
X24339 N24339 N24340 Segment
X24340 N24340 N24341 Segment
X24341 N24341 N24342 Segment
X24342 N24342 N24343 Segment
X24343 N24343 N24344 Segment
X24344 N24344 N24345 Segment
X24345 N24345 N24346 Segment
X24346 N24346 N24347 Segment
X24347 N24347 N24348 Segment
X24348 N24348 N24349 Segment
X24349 N24349 N24350 Segment
X24350 N24350 N24351 Segment
X24351 N24351 N24352 Segment
X24352 N24352 N24353 Segment
X24353 N24353 N24354 Segment
X24354 N24354 N24355 Segment
X24355 N24355 N24356 Segment
X24356 N24356 N24357 Segment
X24357 N24357 N24358 Segment
X24358 N24358 N24359 Segment
X24359 N24359 N24360 Segment
X24360 N24360 N24361 Segment
X24361 N24361 N24362 Segment
X24362 N24362 N24363 Segment
X24363 N24363 N24364 Segment
X24364 N24364 N24365 Segment
X24365 N24365 N24366 Segment
X24366 N24366 N24367 Segment
X24367 N24367 N24368 Segment
X24368 N24368 N24369 Segment
X24369 N24369 N24370 Segment
X24370 N24370 N24371 Segment
X24371 N24371 N24372 Segment
X24372 N24372 N24373 Segment
X24373 N24373 N24374 Segment
X24374 N24374 N24375 Segment
X24375 N24375 N24376 Segment
X24376 N24376 N24377 Segment
X24377 N24377 N24378 Segment
X24378 N24378 N24379 Segment
X24379 N24379 N24380 Segment
X24380 N24380 N24381 Segment
X24381 N24381 N24382 Segment
X24382 N24382 N24383 Segment
X24383 N24383 N24384 Segment
X24384 N24384 N24385 Segment
X24385 N24385 N24386 Segment
X24386 N24386 N24387 Segment
X24387 N24387 N24388 Segment
X24388 N24388 N24389 Segment
X24389 N24389 N24390 Segment
X24390 N24390 N24391 Segment
X24391 N24391 N24392 Segment
X24392 N24392 N24393 Segment
X24393 N24393 N24394 Segment
X24394 N24394 N24395 Segment
X24395 N24395 N24396 Segment
X24396 N24396 N24397 Segment
X24397 N24397 N24398 Segment
X24398 N24398 N24399 Segment
X24399 N24399 N24400 Segment
X24400 N24400 N24401 Segment
X24401 N24401 N24402 Segment
X24402 N24402 N24403 Segment
X24403 N24403 N24404 Segment
X24404 N24404 N24405 Segment
X24405 N24405 N24406 Segment
X24406 N24406 N24407 Segment
X24407 N24407 N24408 Segment
X24408 N24408 N24409 Segment
X24409 N24409 N24410 Segment
X24410 N24410 N24411 Segment
X24411 N24411 N24412 Segment
X24412 N24412 N24413 Segment
X24413 N24413 N24414 Segment
X24414 N24414 N24415 Segment
X24415 N24415 N24416 Segment
X24416 N24416 N24417 Segment
X24417 N24417 N24418 Segment
X24418 N24418 N24419 Segment
X24419 N24419 N24420 Segment
X24420 N24420 N24421 Segment
X24421 N24421 N24422 Segment
X24422 N24422 N24423 Segment
X24423 N24423 N24424 Segment
X24424 N24424 N24425 Segment
X24425 N24425 N24426 Segment
X24426 N24426 N24427 Segment
X24427 N24427 N24428 Segment
X24428 N24428 N24429 Segment
X24429 N24429 N24430 Segment
X24430 N24430 N24431 Segment
X24431 N24431 N24432 Segment
X24432 N24432 N24433 Segment
X24433 N24433 N24434 Segment
X24434 N24434 N24435 Segment
X24435 N24435 N24436 Segment
X24436 N24436 N24437 Segment
X24437 N24437 N24438 Segment
X24438 N24438 N24439 Segment
X24439 N24439 N24440 Segment
X24440 N24440 N24441 Segment
X24441 N24441 N24442 Segment
X24442 N24442 N24443 Segment
X24443 N24443 N24444 Segment
X24444 N24444 N24445 Segment
X24445 N24445 N24446 Segment
X24446 N24446 N24447 Segment
X24447 N24447 N24448 Segment
X24448 N24448 N24449 Segment
X24449 N24449 N24450 Segment
X24450 N24450 N24451 Segment
X24451 N24451 N24452 Segment
X24452 N24452 N24453 Segment
X24453 N24453 N24454 Segment
X24454 N24454 N24455 Segment
X24455 N24455 N24456 Segment
X24456 N24456 N24457 Segment
X24457 N24457 N24458 Segment
X24458 N24458 N24459 Segment
X24459 N24459 N24460 Segment
X24460 N24460 N24461 Segment
X24461 N24461 N24462 Segment
X24462 N24462 N24463 Segment
X24463 N24463 N24464 Segment
X24464 N24464 N24465 Segment
X24465 N24465 N24466 Segment
X24466 N24466 N24467 Segment
X24467 N24467 N24468 Segment
X24468 N24468 N24469 Segment
X24469 N24469 N24470 Segment
X24470 N24470 N24471 Segment
X24471 N24471 N24472 Segment
X24472 N24472 N24473 Segment
X24473 N24473 N24474 Segment
X24474 N24474 N24475 Segment
X24475 N24475 N24476 Segment
X24476 N24476 N24477 Segment
X24477 N24477 N24478 Segment
X24478 N24478 N24479 Segment
X24479 N24479 N24480 Segment
X24480 N24480 N24481 Segment
X24481 N24481 N24482 Segment
X24482 N24482 N24483 Segment
X24483 N24483 N24484 Segment
X24484 N24484 N24485 Segment
X24485 N24485 N24486 Segment
X24486 N24486 N24487 Segment
X24487 N24487 N24488 Segment
X24488 N24488 N24489 Segment
X24489 N24489 N24490 Segment
X24490 N24490 N24491 Segment
X24491 N24491 N24492 Segment
X24492 N24492 N24493 Segment
X24493 N24493 N24494 Segment
X24494 N24494 N24495 Segment
X24495 N24495 N24496 Segment
X24496 N24496 N24497 Segment
X24497 N24497 N24498 Segment
X24498 N24498 N24499 Segment
X24499 N24499 N24500 Segment
X24500 N24500 N24501 Segment
X24501 N24501 N24502 Segment
X24502 N24502 N24503 Segment
X24503 N24503 N24504 Segment
X24504 N24504 N24505 Segment
X24505 N24505 N24506 Segment
X24506 N24506 N24507 Segment
X24507 N24507 N24508 Segment
X24508 N24508 N24509 Segment
X24509 N24509 N24510 Segment
X24510 N24510 N24511 Segment
X24511 N24511 N24512 Segment
X24512 N24512 N24513 Segment
X24513 N24513 N24514 Segment
X24514 N24514 N24515 Segment
X24515 N24515 N24516 Segment
X24516 N24516 N24517 Segment
X24517 N24517 N24518 Segment
X24518 N24518 N24519 Segment
X24519 N24519 N24520 Segment
X24520 N24520 N24521 Segment
X24521 N24521 N24522 Segment
X24522 N24522 N24523 Segment
X24523 N24523 N24524 Segment
X24524 N24524 N24525 Segment
X24525 N24525 N24526 Segment
X24526 N24526 N24527 Segment
X24527 N24527 N24528 Segment
X24528 N24528 N24529 Segment
X24529 N24529 N24530 Segment
X24530 N24530 N24531 Segment
X24531 N24531 N24532 Segment
X24532 N24532 N24533 Segment
X24533 N24533 N24534 Segment
X24534 N24534 N24535 Segment
X24535 N24535 N24536 Segment
X24536 N24536 N24537 Segment
X24537 N24537 N24538 Segment
X24538 N24538 N24539 Segment
X24539 N24539 N24540 Segment
X24540 N24540 N24541 Segment
X24541 N24541 N24542 Segment
X24542 N24542 N24543 Segment
X24543 N24543 N24544 Segment
X24544 N24544 N24545 Segment
X24545 N24545 N24546 Segment
X24546 N24546 N24547 Segment
X24547 N24547 N24548 Segment
X24548 N24548 N24549 Segment
X24549 N24549 N24550 Segment
X24550 N24550 N24551 Segment
X24551 N24551 N24552 Segment
X24552 N24552 N24553 Segment
X24553 N24553 N24554 Segment
X24554 N24554 N24555 Segment
X24555 N24555 N24556 Segment
X24556 N24556 N24557 Segment
X24557 N24557 N24558 Segment
X24558 N24558 N24559 Segment
X24559 N24559 N24560 Segment
X24560 N24560 N24561 Segment
X24561 N24561 N24562 Segment
X24562 N24562 N24563 Segment
X24563 N24563 N24564 Segment
X24564 N24564 N24565 Segment
X24565 N24565 N24566 Segment
X24566 N24566 N24567 Segment
X24567 N24567 N24568 Segment
X24568 N24568 N24569 Segment
X24569 N24569 N24570 Segment
X24570 N24570 N24571 Segment
X24571 N24571 N24572 Segment
X24572 N24572 N24573 Segment
X24573 N24573 N24574 Segment
X24574 N24574 N24575 Segment
X24575 N24575 N24576 Segment
X24576 N24576 N24577 Segment
X24577 N24577 N24578 Segment
X24578 N24578 N24579 Segment
X24579 N24579 N24580 Segment
X24580 N24580 N24581 Segment
X24581 N24581 N24582 Segment
X24582 N24582 N24583 Segment
X24583 N24583 N24584 Segment
X24584 N24584 N24585 Segment
X24585 N24585 N24586 Segment
X24586 N24586 N24587 Segment
X24587 N24587 N24588 Segment
X24588 N24588 N24589 Segment
X24589 N24589 N24590 Segment
X24590 N24590 N24591 Segment
X24591 N24591 N24592 Segment
X24592 N24592 N24593 Segment
X24593 N24593 N24594 Segment
X24594 N24594 N24595 Segment
X24595 N24595 N24596 Segment
X24596 N24596 N24597 Segment
X24597 N24597 N24598 Segment
X24598 N24598 N24599 Segment
X24599 N24599 N24600 Segment
X24600 N24600 N24601 Segment
X24601 N24601 N24602 Segment
X24602 N24602 N24603 Segment
X24603 N24603 N24604 Segment
X24604 N24604 N24605 Segment
X24605 N24605 N24606 Segment
X24606 N24606 N24607 Segment
X24607 N24607 N24608 Segment
X24608 N24608 N24609 Segment
X24609 N24609 N24610 Segment
X24610 N24610 N24611 Segment
X24611 N24611 N24612 Segment
X24612 N24612 N24613 Segment
X24613 N24613 N24614 Segment
X24614 N24614 N24615 Segment
X24615 N24615 N24616 Segment
X24616 N24616 N24617 Segment
X24617 N24617 N24618 Segment
X24618 N24618 N24619 Segment
X24619 N24619 N24620 Segment
X24620 N24620 N24621 Segment
X24621 N24621 N24622 Segment
X24622 N24622 N24623 Segment
X24623 N24623 N24624 Segment
X24624 N24624 N24625 Segment
X24625 N24625 N24626 Segment
X24626 N24626 N24627 Segment
X24627 N24627 N24628 Segment
X24628 N24628 N24629 Segment
X24629 N24629 N24630 Segment
X24630 N24630 N24631 Segment
X24631 N24631 N24632 Segment
X24632 N24632 N24633 Segment
X24633 N24633 N24634 Segment
X24634 N24634 N24635 Segment
X24635 N24635 N24636 Segment
X24636 N24636 N24637 Segment
X24637 N24637 N24638 Segment
X24638 N24638 N24639 Segment
X24639 N24639 N24640 Segment
X24640 N24640 N24641 Segment
X24641 N24641 N24642 Segment
X24642 N24642 N24643 Segment
X24643 N24643 N24644 Segment
X24644 N24644 N24645 Segment
X24645 N24645 N24646 Segment
X24646 N24646 N24647 Segment
X24647 N24647 N24648 Segment
X24648 N24648 N24649 Segment
X24649 N24649 N24650 Segment
X24650 N24650 N24651 Segment
X24651 N24651 N24652 Segment
X24652 N24652 N24653 Segment
X24653 N24653 N24654 Segment
X24654 N24654 N24655 Segment
X24655 N24655 N24656 Segment
X24656 N24656 N24657 Segment
X24657 N24657 N24658 Segment
X24658 N24658 N24659 Segment
X24659 N24659 N24660 Segment
X24660 N24660 N24661 Segment
X24661 N24661 N24662 Segment
X24662 N24662 N24663 Segment
X24663 N24663 N24664 Segment
X24664 N24664 N24665 Segment
X24665 N24665 N24666 Segment
X24666 N24666 N24667 Segment
X24667 N24667 N24668 Segment
X24668 N24668 N24669 Segment
X24669 N24669 N24670 Segment
X24670 N24670 N24671 Segment
X24671 N24671 N24672 Segment
X24672 N24672 N24673 Segment
X24673 N24673 N24674 Segment
X24674 N24674 N24675 Segment
X24675 N24675 N24676 Segment
X24676 N24676 N24677 Segment
X24677 N24677 N24678 Segment
X24678 N24678 N24679 Segment
X24679 N24679 N24680 Segment
X24680 N24680 N24681 Segment
X24681 N24681 N24682 Segment
X24682 N24682 N24683 Segment
X24683 N24683 N24684 Segment
X24684 N24684 N24685 Segment
X24685 N24685 N24686 Segment
X24686 N24686 N24687 Segment
X24687 N24687 N24688 Segment
X24688 N24688 N24689 Segment
X24689 N24689 N24690 Segment
X24690 N24690 N24691 Segment
X24691 N24691 N24692 Segment
X24692 N24692 N24693 Segment
X24693 N24693 N24694 Segment
X24694 N24694 N24695 Segment
X24695 N24695 N24696 Segment
X24696 N24696 N24697 Segment
X24697 N24697 N24698 Segment
X24698 N24698 N24699 Segment
X24699 N24699 N24700 Segment
X24700 N24700 N24701 Segment
X24701 N24701 N24702 Segment
X24702 N24702 N24703 Segment
X24703 N24703 N24704 Segment
X24704 N24704 N24705 Segment
X24705 N24705 N24706 Segment
X24706 N24706 N24707 Segment
X24707 N24707 N24708 Segment
X24708 N24708 N24709 Segment
X24709 N24709 N24710 Segment
X24710 N24710 N24711 Segment
X24711 N24711 N24712 Segment
X24712 N24712 N24713 Segment
X24713 N24713 N24714 Segment
X24714 N24714 N24715 Segment
X24715 N24715 N24716 Segment
X24716 N24716 N24717 Segment
X24717 N24717 N24718 Segment
X24718 N24718 N24719 Segment
X24719 N24719 N24720 Segment
X24720 N24720 N24721 Segment
X24721 N24721 N24722 Segment
X24722 N24722 N24723 Segment
X24723 N24723 N24724 Segment
X24724 N24724 N24725 Segment
X24725 N24725 N24726 Segment
X24726 N24726 N24727 Segment
X24727 N24727 N24728 Segment
X24728 N24728 N24729 Segment
X24729 N24729 N24730 Segment
X24730 N24730 N24731 Segment
X24731 N24731 N24732 Segment
X24732 N24732 N24733 Segment
X24733 N24733 N24734 Segment
X24734 N24734 N24735 Segment
X24735 N24735 N24736 Segment
X24736 N24736 N24737 Segment
X24737 N24737 N24738 Segment
X24738 N24738 N24739 Segment
X24739 N24739 N24740 Segment
X24740 N24740 N24741 Segment
X24741 N24741 N24742 Segment
X24742 N24742 N24743 Segment
X24743 N24743 N24744 Segment
X24744 N24744 N24745 Segment
X24745 N24745 N24746 Segment
X24746 N24746 N24747 Segment
X24747 N24747 N24748 Segment
X24748 N24748 N24749 Segment
X24749 N24749 N24750 Segment
X24750 N24750 N24751 Segment
X24751 N24751 N24752 Segment
X24752 N24752 N24753 Segment
X24753 N24753 N24754 Segment
X24754 N24754 N24755 Segment
X24755 N24755 N24756 Segment
X24756 N24756 N24757 Segment
X24757 N24757 N24758 Segment
X24758 N24758 N24759 Segment
X24759 N24759 N24760 Segment
X24760 N24760 N24761 Segment
X24761 N24761 N24762 Segment
X24762 N24762 N24763 Segment
X24763 N24763 N24764 Segment
X24764 N24764 N24765 Segment
X24765 N24765 N24766 Segment
X24766 N24766 N24767 Segment
X24767 N24767 N24768 Segment
X24768 N24768 N24769 Segment
X24769 N24769 N24770 Segment
X24770 N24770 N24771 Segment
X24771 N24771 N24772 Segment
X24772 N24772 N24773 Segment
X24773 N24773 N24774 Segment
X24774 N24774 N24775 Segment
X24775 N24775 N24776 Segment
X24776 N24776 N24777 Segment
X24777 N24777 N24778 Segment
X24778 N24778 N24779 Segment
X24779 N24779 N24780 Segment
X24780 N24780 N24781 Segment
X24781 N24781 N24782 Segment
X24782 N24782 N24783 Segment
X24783 N24783 N24784 Segment
X24784 N24784 N24785 Segment
X24785 N24785 N24786 Segment
X24786 N24786 N24787 Segment
X24787 N24787 N24788 Segment
X24788 N24788 N24789 Segment
X24789 N24789 N24790 Segment
X24790 N24790 N24791 Segment
X24791 N24791 N24792 Segment
X24792 N24792 N24793 Segment
X24793 N24793 N24794 Segment
X24794 N24794 N24795 Segment
X24795 N24795 N24796 Segment
X24796 N24796 N24797 Segment
X24797 N24797 N24798 Segment
X24798 N24798 N24799 Segment
X24799 N24799 N24800 Segment
X24800 N24800 N24801 Segment
X24801 N24801 N24802 Segment
X24802 N24802 N24803 Segment
X24803 N24803 N24804 Segment
X24804 N24804 N24805 Segment
X24805 N24805 N24806 Segment
X24806 N24806 N24807 Segment
X24807 N24807 N24808 Segment
X24808 N24808 N24809 Segment
X24809 N24809 N24810 Segment
X24810 N24810 N24811 Segment
X24811 N24811 N24812 Segment
X24812 N24812 N24813 Segment
X24813 N24813 N24814 Segment
X24814 N24814 N24815 Segment
X24815 N24815 N24816 Segment
X24816 N24816 N24817 Segment
X24817 N24817 N24818 Segment
X24818 N24818 N24819 Segment
X24819 N24819 N24820 Segment
X24820 N24820 N24821 Segment
X24821 N24821 N24822 Segment
X24822 N24822 N24823 Segment
X24823 N24823 N24824 Segment
X24824 N24824 N24825 Segment
X24825 N24825 N24826 Segment
X24826 N24826 N24827 Segment
X24827 N24827 N24828 Segment
X24828 N24828 N24829 Segment
X24829 N24829 N24830 Segment
X24830 N24830 N24831 Segment
X24831 N24831 N24832 Segment
X24832 N24832 N24833 Segment
X24833 N24833 N24834 Segment
X24834 N24834 N24835 Segment
X24835 N24835 N24836 Segment
X24836 N24836 N24837 Segment
X24837 N24837 N24838 Segment
X24838 N24838 N24839 Segment
X24839 N24839 N24840 Segment
X24840 N24840 N24841 Segment
X24841 N24841 N24842 Segment
X24842 N24842 N24843 Segment
X24843 N24843 N24844 Segment
X24844 N24844 N24845 Segment
X24845 N24845 N24846 Segment
X24846 N24846 N24847 Segment
X24847 N24847 N24848 Segment
X24848 N24848 N24849 Segment
X24849 N24849 N24850 Segment
X24850 N24850 N24851 Segment
X24851 N24851 N24852 Segment
X24852 N24852 N24853 Segment
X24853 N24853 N24854 Segment
X24854 N24854 N24855 Segment
X24855 N24855 N24856 Segment
X24856 N24856 N24857 Segment
X24857 N24857 N24858 Segment
X24858 N24858 N24859 Segment
X24859 N24859 N24860 Segment
X24860 N24860 N24861 Segment
X24861 N24861 N24862 Segment
X24862 N24862 N24863 Segment
X24863 N24863 N24864 Segment
X24864 N24864 N24865 Segment
X24865 N24865 N24866 Segment
X24866 N24866 N24867 Segment
X24867 N24867 N24868 Segment
X24868 N24868 N24869 Segment
X24869 N24869 N24870 Segment
X24870 N24870 N24871 Segment
X24871 N24871 N24872 Segment
X24872 N24872 N24873 Segment
X24873 N24873 N24874 Segment
X24874 N24874 N24875 Segment
X24875 N24875 N24876 Segment
X24876 N24876 N24877 Segment
X24877 N24877 N24878 Segment
X24878 N24878 N24879 Segment
X24879 N24879 N24880 Segment
X24880 N24880 N24881 Segment
X24881 N24881 N24882 Segment
X24882 N24882 N24883 Segment
X24883 N24883 N24884 Segment
X24884 N24884 N24885 Segment
X24885 N24885 N24886 Segment
X24886 N24886 N24887 Segment
X24887 N24887 N24888 Segment
X24888 N24888 N24889 Segment
X24889 N24889 N24890 Segment
X24890 N24890 N24891 Segment
X24891 N24891 N24892 Segment
X24892 N24892 N24893 Segment
X24893 N24893 N24894 Segment
X24894 N24894 N24895 Segment
X24895 N24895 N24896 Segment
X24896 N24896 N24897 Segment
X24897 N24897 N24898 Segment
X24898 N24898 N24899 Segment
X24899 N24899 N24900 Segment
X24900 N24900 N24901 Segment
X24901 N24901 N24902 Segment
X24902 N24902 N24903 Segment
X24903 N24903 N24904 Segment
X24904 N24904 N24905 Segment
X24905 N24905 N24906 Segment
X24906 N24906 N24907 Segment
X24907 N24907 N24908 Segment
X24908 N24908 N24909 Segment
X24909 N24909 N24910 Segment
X24910 N24910 N24911 Segment
X24911 N24911 N24912 Segment
X24912 N24912 N24913 Segment
X24913 N24913 N24914 Segment
X24914 N24914 N24915 Segment
X24915 N24915 N24916 Segment
X24916 N24916 N24917 Segment
X24917 N24917 N24918 Segment
X24918 N24918 N24919 Segment
X24919 N24919 N24920 Segment
X24920 N24920 N24921 Segment
X24921 N24921 N24922 Segment
X24922 N24922 N24923 Segment
X24923 N24923 N24924 Segment
X24924 N24924 N24925 Segment
X24925 N24925 N24926 Segment
X24926 N24926 N24927 Segment
X24927 N24927 N24928 Segment
X24928 N24928 N24929 Segment
X24929 N24929 N24930 Segment
X24930 N24930 N24931 Segment
X24931 N24931 N24932 Segment
X24932 N24932 N24933 Segment
X24933 N24933 N24934 Segment
X24934 N24934 N24935 Segment
X24935 N24935 N24936 Segment
X24936 N24936 N24937 Segment
X24937 N24937 N24938 Segment
X24938 N24938 N24939 Segment
X24939 N24939 N24940 Segment
X24940 N24940 N24941 Segment
X24941 N24941 N24942 Segment
X24942 N24942 N24943 Segment
X24943 N24943 N24944 Segment
X24944 N24944 N24945 Segment
X24945 N24945 N24946 Segment
X24946 N24946 N24947 Segment
X24947 N24947 N24948 Segment
X24948 N24948 N24949 Segment
X24949 N24949 N24950 Segment
X24950 N24950 N24951 Segment
X24951 N24951 N24952 Segment
X24952 N24952 N24953 Segment
X24953 N24953 N24954 Segment
X24954 N24954 N24955 Segment
X24955 N24955 N24956 Segment
X24956 N24956 N24957 Segment
X24957 N24957 N24958 Segment
X24958 N24958 N24959 Segment
X24959 N24959 N24960 Segment
X24960 N24960 N24961 Segment
X24961 N24961 N24962 Segment
X24962 N24962 N24963 Segment
X24963 N24963 N24964 Segment
X24964 N24964 N24965 Segment
X24965 N24965 N24966 Segment
X24966 N24966 N24967 Segment
X24967 N24967 N24968 Segment
X24968 N24968 N24969 Segment
X24969 N24969 N24970 Segment
X24970 N24970 N24971 Segment
X24971 N24971 N24972 Segment
X24972 N24972 N24973 Segment
X24973 N24973 N24974 Segment
X24974 N24974 N24975 Segment
X24975 N24975 N24976 Segment
X24976 N24976 N24977 Segment
X24977 N24977 N24978 Segment
X24978 N24978 N24979 Segment
X24979 N24979 N24980 Segment
X24980 N24980 N24981 Segment
X24981 N24981 N24982 Segment
X24982 N24982 N24983 Segment
X24983 N24983 N24984 Segment
X24984 N24984 N24985 Segment
X24985 N24985 N24986 Segment
X24986 N24986 N24987 Segment
X24987 N24987 N24988 Segment
X24988 N24988 N24989 Segment
X24989 N24989 N24990 Segment
X24990 N24990 N24991 Segment
X24991 N24991 N24992 Segment
X24992 N24992 N24993 Segment
X24993 N24993 N24994 Segment
X24994 N24994 N24995 Segment
X24995 N24995 N24996 Segment
X24996 N24996 N24997 Segment
X24997 N24997 N24998 Segment
X24998 N24998 N24999 Segment
X24999 N24999 N25000 Segment
X25000 N25000 N25001 Segment
X25001 N25001 N25002 Segment
X25002 N25002 N25003 Segment
X25003 N25003 N25004 Segment
X25004 N25004 N25005 Segment
X25005 N25005 N25006 Segment
X25006 N25006 N25007 Segment
X25007 N25007 N25008 Segment
X25008 N25008 N25009 Segment
X25009 N25009 N25010 Segment
X25010 N25010 N25011 Segment
X25011 N25011 N25012 Segment
X25012 N25012 N25013 Segment
X25013 N25013 N25014 Segment
X25014 N25014 N25015 Segment
X25015 N25015 N25016 Segment
X25016 N25016 N25017 Segment
X25017 N25017 N25018 Segment
X25018 N25018 N25019 Segment
X25019 N25019 N25020 Segment
X25020 N25020 N25021 Segment
X25021 N25021 N25022 Segment
X25022 N25022 N25023 Segment
X25023 N25023 N25024 Segment
X25024 N25024 N25025 Segment
X25025 N25025 N25026 Segment
X25026 N25026 N25027 Segment
X25027 N25027 N25028 Segment
X25028 N25028 N25029 Segment
X25029 N25029 N25030 Segment
X25030 N25030 N25031 Segment
X25031 N25031 N25032 Segment
X25032 N25032 N25033 Segment
X25033 N25033 N25034 Segment
X25034 N25034 N25035 Segment
X25035 N25035 N25036 Segment
X25036 N25036 N25037 Segment
X25037 N25037 N25038 Segment
X25038 N25038 N25039 Segment
X25039 N25039 N25040 Segment
X25040 N25040 N25041 Segment
X25041 N25041 N25042 Segment
X25042 N25042 N25043 Segment
X25043 N25043 N25044 Segment
X25044 N25044 N25045 Segment
X25045 N25045 N25046 Segment
X25046 N25046 N25047 Segment
X25047 N25047 N25048 Segment
X25048 N25048 N25049 Segment
X25049 N25049 N25050 Segment
X25050 N25050 N25051 Segment
X25051 N25051 N25052 Segment
X25052 N25052 N25053 Segment
X25053 N25053 N25054 Segment
X25054 N25054 N25055 Segment
X25055 N25055 N25056 Segment
X25056 N25056 N25057 Segment
X25057 N25057 N25058 Segment
X25058 N25058 N25059 Segment
X25059 N25059 N25060 Segment
X25060 N25060 N25061 Segment
X25061 N25061 N25062 Segment
X25062 N25062 N25063 Segment
X25063 N25063 N25064 Segment
X25064 N25064 N25065 Segment
X25065 N25065 N25066 Segment
X25066 N25066 N25067 Segment
X25067 N25067 N25068 Segment
X25068 N25068 N25069 Segment
X25069 N25069 N25070 Segment
X25070 N25070 N25071 Segment
X25071 N25071 N25072 Segment
X25072 N25072 N25073 Segment
X25073 N25073 N25074 Segment
X25074 N25074 N25075 Segment
X25075 N25075 N25076 Segment
X25076 N25076 N25077 Segment
X25077 N25077 N25078 Segment
X25078 N25078 N25079 Segment
X25079 N25079 N25080 Segment
X25080 N25080 N25081 Segment
X25081 N25081 N25082 Segment
X25082 N25082 N25083 Segment
X25083 N25083 N25084 Segment
X25084 N25084 N25085 Segment
X25085 N25085 N25086 Segment
X25086 N25086 N25087 Segment
X25087 N25087 N25088 Segment
X25088 N25088 N25089 Segment
X25089 N25089 N25090 Segment
X25090 N25090 N25091 Segment
X25091 N25091 N25092 Segment
X25092 N25092 N25093 Segment
X25093 N25093 N25094 Segment
X25094 N25094 N25095 Segment
X25095 N25095 N25096 Segment
X25096 N25096 N25097 Segment
X25097 N25097 N25098 Segment
X25098 N25098 N25099 Segment
X25099 N25099 N25100 Segment
X25100 N25100 N25101 Segment
X25101 N25101 N25102 Segment
X25102 N25102 N25103 Segment
X25103 N25103 N25104 Segment
X25104 N25104 N25105 Segment
X25105 N25105 N25106 Segment
X25106 N25106 N25107 Segment
X25107 N25107 N25108 Segment
X25108 N25108 N25109 Segment
X25109 N25109 N25110 Segment
X25110 N25110 N25111 Segment
X25111 N25111 N25112 Segment
X25112 N25112 N25113 Segment
X25113 N25113 N25114 Segment
X25114 N25114 N25115 Segment
X25115 N25115 N25116 Segment
X25116 N25116 N25117 Segment
X25117 N25117 N25118 Segment
X25118 N25118 N25119 Segment
X25119 N25119 N25120 Segment
X25120 N25120 N25121 Segment
X25121 N25121 N25122 Segment
X25122 N25122 N25123 Segment
X25123 N25123 N25124 Segment
X25124 N25124 N25125 Segment
X25125 N25125 N25126 Segment
X25126 N25126 N25127 Segment
X25127 N25127 N25128 Segment
X25128 N25128 N25129 Segment
X25129 N25129 N25130 Segment
X25130 N25130 N25131 Segment
X25131 N25131 N25132 Segment
X25132 N25132 N25133 Segment
X25133 N25133 N25134 Segment
X25134 N25134 N25135 Segment
X25135 N25135 N25136 Segment
X25136 N25136 N25137 Segment
X25137 N25137 N25138 Segment
X25138 N25138 N25139 Segment
X25139 N25139 N25140 Segment
X25140 N25140 N25141 Segment
X25141 N25141 N25142 Segment
X25142 N25142 N25143 Segment
X25143 N25143 N25144 Segment
X25144 N25144 N25145 Segment
X25145 N25145 N25146 Segment
X25146 N25146 N25147 Segment
X25147 N25147 N25148 Segment
X25148 N25148 N25149 Segment
X25149 N25149 N25150 Segment
X25150 N25150 N25151 Segment
X25151 N25151 N25152 Segment
X25152 N25152 N25153 Segment
X25153 N25153 N25154 Segment
X25154 N25154 N25155 Segment
X25155 N25155 N25156 Segment
X25156 N25156 N25157 Segment
X25157 N25157 N25158 Segment
X25158 N25158 N25159 Segment
X25159 N25159 N25160 Segment
X25160 N25160 N25161 Segment
X25161 N25161 N25162 Segment
X25162 N25162 N25163 Segment
X25163 N25163 N25164 Segment
X25164 N25164 N25165 Segment
X25165 N25165 N25166 Segment
X25166 N25166 N25167 Segment
X25167 N25167 N25168 Segment
X25168 N25168 N25169 Segment
X25169 N25169 N25170 Segment
X25170 N25170 N25171 Segment
X25171 N25171 N25172 Segment
X25172 N25172 N25173 Segment
X25173 N25173 N25174 Segment
X25174 N25174 N25175 Segment
X25175 N25175 N25176 Segment
X25176 N25176 N25177 Segment
X25177 N25177 N25178 Segment
X25178 N25178 N25179 Segment
X25179 N25179 N25180 Segment
X25180 N25180 N25181 Segment
X25181 N25181 N25182 Segment
X25182 N25182 N25183 Segment
X25183 N25183 N25184 Segment
X25184 N25184 N25185 Segment
X25185 N25185 N25186 Segment
X25186 N25186 N25187 Segment
X25187 N25187 N25188 Segment
X25188 N25188 N25189 Segment
X25189 N25189 N25190 Segment
X25190 N25190 N25191 Segment
X25191 N25191 N25192 Segment
X25192 N25192 N25193 Segment
X25193 N25193 N25194 Segment
X25194 N25194 N25195 Segment
X25195 N25195 N25196 Segment
X25196 N25196 N25197 Segment
X25197 N25197 N25198 Segment
X25198 N25198 N25199 Segment
X25199 N25199 N25200 Segment
X25200 N25200 N25201 Segment
X25201 N25201 N25202 Segment
X25202 N25202 N25203 Segment
X25203 N25203 N25204 Segment
X25204 N25204 N25205 Segment
X25205 N25205 N25206 Segment
X25206 N25206 N25207 Segment
X25207 N25207 N25208 Segment
X25208 N25208 N25209 Segment
X25209 N25209 N25210 Segment
X25210 N25210 N25211 Segment
X25211 N25211 N25212 Segment
X25212 N25212 N25213 Segment
X25213 N25213 N25214 Segment
X25214 N25214 N25215 Segment
X25215 N25215 N25216 Segment
X25216 N25216 N25217 Segment
X25217 N25217 N25218 Segment
X25218 N25218 N25219 Segment
X25219 N25219 N25220 Segment
X25220 N25220 N25221 Segment
X25221 N25221 N25222 Segment
X25222 N25222 N25223 Segment
X25223 N25223 N25224 Segment
X25224 N25224 N25225 Segment
X25225 N25225 N25226 Segment
X25226 N25226 N25227 Segment
X25227 N25227 N25228 Segment
X25228 N25228 N25229 Segment
X25229 N25229 N25230 Segment
X25230 N25230 N25231 Segment
X25231 N25231 N25232 Segment
X25232 N25232 N25233 Segment
X25233 N25233 N25234 Segment
X25234 N25234 N25235 Segment
X25235 N25235 N25236 Segment
X25236 N25236 N25237 Segment
X25237 N25237 N25238 Segment
X25238 N25238 N25239 Segment
X25239 N25239 N25240 Segment
X25240 N25240 N25241 Segment
X25241 N25241 N25242 Segment
X25242 N25242 N25243 Segment
X25243 N25243 N25244 Segment
X25244 N25244 N25245 Segment
X25245 N25245 N25246 Segment
X25246 N25246 N25247 Segment
X25247 N25247 N25248 Segment
X25248 N25248 N25249 Segment
X25249 N25249 N25250 Segment
X25250 N25250 N25251 Segment
X25251 N25251 N25252 Segment
X25252 N25252 N25253 Segment
X25253 N25253 N25254 Segment
X25254 N25254 N25255 Segment
X25255 N25255 N25256 Segment
X25256 N25256 N25257 Segment
X25257 N25257 N25258 Segment
X25258 N25258 N25259 Segment
X25259 N25259 N25260 Segment
X25260 N25260 N25261 Segment
X25261 N25261 N25262 Segment
X25262 N25262 N25263 Segment
X25263 N25263 N25264 Segment
X25264 N25264 N25265 Segment
X25265 N25265 N25266 Segment
X25266 N25266 N25267 Segment
X25267 N25267 N25268 Segment
X25268 N25268 N25269 Segment
X25269 N25269 N25270 Segment
X25270 N25270 N25271 Segment
X25271 N25271 N25272 Segment
X25272 N25272 N25273 Segment
X25273 N25273 N25274 Segment
X25274 N25274 N25275 Segment
X25275 N25275 N25276 Segment
X25276 N25276 N25277 Segment
X25277 N25277 N25278 Segment
X25278 N25278 N25279 Segment
X25279 N25279 N25280 Segment
X25280 N25280 N25281 Segment
X25281 N25281 N25282 Segment
X25282 N25282 N25283 Segment
X25283 N25283 N25284 Segment
X25284 N25284 N25285 Segment
X25285 N25285 N25286 Segment
X25286 N25286 N25287 Segment
X25287 N25287 N25288 Segment
X25288 N25288 N25289 Segment
X25289 N25289 N25290 Segment
X25290 N25290 N25291 Segment
X25291 N25291 N25292 Segment
X25292 N25292 N25293 Segment
X25293 N25293 N25294 Segment
X25294 N25294 N25295 Segment
X25295 N25295 N25296 Segment
X25296 N25296 N25297 Segment
X25297 N25297 N25298 Segment
X25298 N25298 N25299 Segment
X25299 N25299 N25300 Segment
X25300 N25300 N25301 Segment
X25301 N25301 N25302 Segment
X25302 N25302 N25303 Segment
X25303 N25303 N25304 Segment
X25304 N25304 N25305 Segment
X25305 N25305 N25306 Segment
X25306 N25306 N25307 Segment
X25307 N25307 N25308 Segment
X25308 N25308 N25309 Segment
X25309 N25309 N25310 Segment
X25310 N25310 N25311 Segment
X25311 N25311 N25312 Segment
X25312 N25312 N25313 Segment
X25313 N25313 N25314 Segment
X25314 N25314 N25315 Segment
X25315 N25315 N25316 Segment
X25316 N25316 N25317 Segment
X25317 N25317 N25318 Segment
X25318 N25318 N25319 Segment
X25319 N25319 N25320 Segment
X25320 N25320 N25321 Segment
X25321 N25321 N25322 Segment
X25322 N25322 N25323 Segment
X25323 N25323 N25324 Segment
X25324 N25324 N25325 Segment
X25325 N25325 N25326 Segment
X25326 N25326 N25327 Segment
X25327 N25327 N25328 Segment
X25328 N25328 N25329 Segment
X25329 N25329 N25330 Segment
X25330 N25330 N25331 Segment
X25331 N25331 N25332 Segment
X25332 N25332 N25333 Segment
X25333 N25333 N25334 Segment
X25334 N25334 N25335 Segment
X25335 N25335 N25336 Segment
X25336 N25336 N25337 Segment
X25337 N25337 N25338 Segment
X25338 N25338 N25339 Segment
X25339 N25339 N25340 Segment
X25340 N25340 N25341 Segment
X25341 N25341 N25342 Segment
X25342 N25342 N25343 Segment
X25343 N25343 N25344 Segment
X25344 N25344 N25345 Segment
X25345 N25345 N25346 Segment
X25346 N25346 N25347 Segment
X25347 N25347 N25348 Segment
X25348 N25348 N25349 Segment
X25349 N25349 N25350 Segment
X25350 N25350 N25351 Segment
X25351 N25351 N25352 Segment
X25352 N25352 N25353 Segment
X25353 N25353 N25354 Segment
X25354 N25354 N25355 Segment
X25355 N25355 N25356 Segment
X25356 N25356 N25357 Segment
X25357 N25357 N25358 Segment
X25358 N25358 N25359 Segment
X25359 N25359 N25360 Segment
X25360 N25360 N25361 Segment
X25361 N25361 N25362 Segment
X25362 N25362 N25363 Segment
X25363 N25363 N25364 Segment
X25364 N25364 N25365 Segment
X25365 N25365 N25366 Segment
X25366 N25366 N25367 Segment
X25367 N25367 N25368 Segment
X25368 N25368 N25369 Segment
X25369 N25369 N25370 Segment
X25370 N25370 N25371 Segment
X25371 N25371 N25372 Segment
X25372 N25372 N25373 Segment
X25373 N25373 N25374 Segment
X25374 N25374 N25375 Segment
X25375 N25375 N25376 Segment
X25376 N25376 N25377 Segment
X25377 N25377 N25378 Segment
X25378 N25378 N25379 Segment
X25379 N25379 N25380 Segment
X25380 N25380 N25381 Segment
X25381 N25381 N25382 Segment
X25382 N25382 N25383 Segment
X25383 N25383 N25384 Segment
X25384 N25384 N25385 Segment
X25385 N25385 N25386 Segment
X25386 N25386 N25387 Segment
X25387 N25387 N25388 Segment
X25388 N25388 N25389 Segment
X25389 N25389 N25390 Segment
X25390 N25390 N25391 Segment
X25391 N25391 N25392 Segment
X25392 N25392 N25393 Segment
X25393 N25393 N25394 Segment
X25394 N25394 N25395 Segment
X25395 N25395 N25396 Segment
X25396 N25396 N25397 Segment
X25397 N25397 N25398 Segment
X25398 N25398 N25399 Segment
X25399 N25399 N25400 Segment
X25400 N25400 N25401 Segment
X25401 N25401 N25402 Segment
X25402 N25402 N25403 Segment
X25403 N25403 N25404 Segment
X25404 N25404 N25405 Segment
X25405 N25405 N25406 Segment
X25406 N25406 N25407 Segment
X25407 N25407 N25408 Segment
X25408 N25408 N25409 Segment
X25409 N25409 N25410 Segment
X25410 N25410 N25411 Segment
X25411 N25411 N25412 Segment
X25412 N25412 N25413 Segment
X25413 N25413 N25414 Segment
X25414 N25414 N25415 Segment
X25415 N25415 N25416 Segment
X25416 N25416 N25417 Segment
X25417 N25417 N25418 Segment
X25418 N25418 N25419 Segment
X25419 N25419 N25420 Segment
X25420 N25420 N25421 Segment
X25421 N25421 N25422 Segment
X25422 N25422 N25423 Segment
X25423 N25423 N25424 Segment
X25424 N25424 N25425 Segment
X25425 N25425 N25426 Segment
X25426 N25426 N25427 Segment
X25427 N25427 N25428 Segment
X25428 N25428 N25429 Segment
X25429 N25429 N25430 Segment
X25430 N25430 N25431 Segment
X25431 N25431 N25432 Segment
X25432 N25432 N25433 Segment
X25433 N25433 N25434 Segment
X25434 N25434 N25435 Segment
X25435 N25435 N25436 Segment
X25436 N25436 N25437 Segment
X25437 N25437 N25438 Segment
X25438 N25438 N25439 Segment
X25439 N25439 N25440 Segment
X25440 N25440 N25441 Segment
X25441 N25441 N25442 Segment
X25442 N25442 N25443 Segment
X25443 N25443 N25444 Segment
X25444 N25444 N25445 Segment
X25445 N25445 N25446 Segment
X25446 N25446 N25447 Segment
X25447 N25447 N25448 Segment
X25448 N25448 N25449 Segment
X25449 N25449 N25450 Segment
X25450 N25450 N25451 Segment
X25451 N25451 N25452 Segment
X25452 N25452 N25453 Segment
X25453 N25453 N25454 Segment
X25454 N25454 N25455 Segment
X25455 N25455 N25456 Segment
X25456 N25456 N25457 Segment
X25457 N25457 N25458 Segment
X25458 N25458 N25459 Segment
X25459 N25459 N25460 Segment
X25460 N25460 N25461 Segment
X25461 N25461 N25462 Segment
X25462 N25462 N25463 Segment
X25463 N25463 N25464 Segment
X25464 N25464 N25465 Segment
X25465 N25465 N25466 Segment
X25466 N25466 N25467 Segment
X25467 N25467 N25468 Segment
X25468 N25468 N25469 Segment
X25469 N25469 N25470 Segment
X25470 N25470 N25471 Segment
X25471 N25471 N25472 Segment
X25472 N25472 N25473 Segment
X25473 N25473 N25474 Segment
X25474 N25474 N25475 Segment
X25475 N25475 N25476 Segment
X25476 N25476 N25477 Segment
X25477 N25477 N25478 Segment
X25478 N25478 N25479 Segment
X25479 N25479 N25480 Segment
X25480 N25480 N25481 Segment
X25481 N25481 N25482 Segment
X25482 N25482 N25483 Segment
X25483 N25483 N25484 Segment
X25484 N25484 N25485 Segment
X25485 N25485 N25486 Segment
X25486 N25486 N25487 Segment
X25487 N25487 N25488 Segment
X25488 N25488 N25489 Segment
X25489 N25489 N25490 Segment
X25490 N25490 N25491 Segment
X25491 N25491 N25492 Segment
X25492 N25492 N25493 Segment
X25493 N25493 N25494 Segment
X25494 N25494 N25495 Segment
X25495 N25495 N25496 Segment
X25496 N25496 N25497 Segment
X25497 N25497 N25498 Segment
X25498 N25498 N25499 Segment
X25499 N25499 N25500 Segment
X25500 N25500 N25501 Segment
X25501 N25501 N25502 Segment
X25502 N25502 N25503 Segment
X25503 N25503 N25504 Segment
X25504 N25504 N25505 Segment
X25505 N25505 N25506 Segment
X25506 N25506 N25507 Segment
X25507 N25507 N25508 Segment
X25508 N25508 N25509 Segment
X25509 N25509 N25510 Segment
X25510 N25510 N25511 Segment
X25511 N25511 N25512 Segment
X25512 N25512 N25513 Segment
X25513 N25513 N25514 Segment
X25514 N25514 N25515 Segment
X25515 N25515 N25516 Segment
X25516 N25516 N25517 Segment
X25517 N25517 N25518 Segment
X25518 N25518 N25519 Segment
X25519 N25519 N25520 Segment
X25520 N25520 N25521 Segment
X25521 N25521 N25522 Segment
X25522 N25522 N25523 Segment
X25523 N25523 N25524 Segment
X25524 N25524 N25525 Segment
X25525 N25525 N25526 Segment
X25526 N25526 N25527 Segment
X25527 N25527 N25528 Segment
X25528 N25528 N25529 Segment
X25529 N25529 N25530 Segment
X25530 N25530 N25531 Segment
X25531 N25531 N25532 Segment
X25532 N25532 N25533 Segment
X25533 N25533 N25534 Segment
X25534 N25534 N25535 Segment
X25535 N25535 N25536 Segment
X25536 N25536 N25537 Segment
X25537 N25537 N25538 Segment
X25538 N25538 N25539 Segment
X25539 N25539 N25540 Segment
X25540 N25540 N25541 Segment
X25541 N25541 N25542 Segment
X25542 N25542 N25543 Segment
X25543 N25543 N25544 Segment
X25544 N25544 N25545 Segment
X25545 N25545 N25546 Segment
X25546 N25546 N25547 Segment
X25547 N25547 N25548 Segment
X25548 N25548 N25549 Segment
X25549 N25549 N25550 Segment
X25550 N25550 N25551 Segment
X25551 N25551 N25552 Segment
X25552 N25552 N25553 Segment
X25553 N25553 N25554 Segment
X25554 N25554 N25555 Segment
X25555 N25555 N25556 Segment
X25556 N25556 N25557 Segment
X25557 N25557 N25558 Segment
X25558 N25558 N25559 Segment
X25559 N25559 N25560 Segment
X25560 N25560 N25561 Segment
X25561 N25561 N25562 Segment
X25562 N25562 N25563 Segment
X25563 N25563 N25564 Segment
X25564 N25564 N25565 Segment
X25565 N25565 N25566 Segment
X25566 N25566 N25567 Segment
X25567 N25567 N25568 Segment
X25568 N25568 N25569 Segment
X25569 N25569 N25570 Segment
X25570 N25570 N25571 Segment
X25571 N25571 N25572 Segment
X25572 N25572 N25573 Segment
X25573 N25573 N25574 Segment
X25574 N25574 N25575 Segment
X25575 N25575 N25576 Segment
X25576 N25576 N25577 Segment
X25577 N25577 N25578 Segment
X25578 N25578 N25579 Segment
X25579 N25579 N25580 Segment
X25580 N25580 N25581 Segment
X25581 N25581 N25582 Segment
X25582 N25582 N25583 Segment
X25583 N25583 N25584 Segment
X25584 N25584 N25585 Segment
X25585 N25585 N25586 Segment
X25586 N25586 N25587 Segment
X25587 N25587 N25588 Segment
X25588 N25588 N25589 Segment
X25589 N25589 N25590 Segment
X25590 N25590 N25591 Segment
X25591 N25591 N25592 Segment
X25592 N25592 N25593 Segment
X25593 N25593 N25594 Segment
X25594 N25594 N25595 Segment
X25595 N25595 N25596 Segment
X25596 N25596 N25597 Segment
X25597 N25597 N25598 Segment
X25598 N25598 N25599 Segment
X25599 N25599 N25600 Segment
X25600 N25600 N25601 Segment
X25601 N25601 N25602 Segment
X25602 N25602 N25603 Segment
X25603 N25603 N25604 Segment
X25604 N25604 N25605 Segment
X25605 N25605 N25606 Segment
X25606 N25606 N25607 Segment
X25607 N25607 N25608 Segment
X25608 N25608 N25609 Segment
X25609 N25609 N25610 Segment
X25610 N25610 N25611 Segment
X25611 N25611 N25612 Segment
X25612 N25612 N25613 Segment
X25613 N25613 N25614 Segment
X25614 N25614 N25615 Segment
X25615 N25615 N25616 Segment
X25616 N25616 N25617 Segment
X25617 N25617 N25618 Segment
X25618 N25618 N25619 Segment
X25619 N25619 N25620 Segment
X25620 N25620 N25621 Segment
X25621 N25621 N25622 Segment
X25622 N25622 N25623 Segment
X25623 N25623 N25624 Segment
X25624 N25624 N25625 Segment
X25625 N25625 N25626 Segment
X25626 N25626 N25627 Segment
X25627 N25627 N25628 Segment
X25628 N25628 N25629 Segment
X25629 N25629 N25630 Segment
X25630 N25630 N25631 Segment
X25631 N25631 N25632 Segment
X25632 N25632 N25633 Segment
X25633 N25633 N25634 Segment
X25634 N25634 N25635 Segment
X25635 N25635 N25636 Segment
X25636 N25636 N25637 Segment
X25637 N25637 N25638 Segment
X25638 N25638 N25639 Segment
X25639 N25639 N25640 Segment
X25640 N25640 N25641 Segment
X25641 N25641 N25642 Segment
X25642 N25642 N25643 Segment
X25643 N25643 N25644 Segment
X25644 N25644 N25645 Segment
X25645 N25645 N25646 Segment
X25646 N25646 N25647 Segment
X25647 N25647 N25648 Segment
X25648 N25648 N25649 Segment
X25649 N25649 N25650 Segment
X25650 N25650 N25651 Segment
X25651 N25651 N25652 Segment
X25652 N25652 N25653 Segment
X25653 N25653 N25654 Segment
X25654 N25654 N25655 Segment
X25655 N25655 N25656 Segment
X25656 N25656 N25657 Segment
X25657 N25657 N25658 Segment
X25658 N25658 N25659 Segment
X25659 N25659 N25660 Segment
X25660 N25660 N25661 Segment
X25661 N25661 N25662 Segment
X25662 N25662 N25663 Segment
X25663 N25663 N25664 Segment
X25664 N25664 N25665 Segment
X25665 N25665 N25666 Segment
X25666 N25666 N25667 Segment
X25667 N25667 N25668 Segment
X25668 N25668 N25669 Segment
X25669 N25669 N25670 Segment
X25670 N25670 N25671 Segment
X25671 N25671 N25672 Segment
X25672 N25672 N25673 Segment
X25673 N25673 N25674 Segment
X25674 N25674 N25675 Segment
X25675 N25675 N25676 Segment
X25676 N25676 N25677 Segment
X25677 N25677 N25678 Segment
X25678 N25678 N25679 Segment
X25679 N25679 N25680 Segment
X25680 N25680 N25681 Segment
X25681 N25681 N25682 Segment
X25682 N25682 N25683 Segment
X25683 N25683 N25684 Segment
X25684 N25684 N25685 Segment
X25685 N25685 N25686 Segment
X25686 N25686 N25687 Segment
X25687 N25687 N25688 Segment
X25688 N25688 N25689 Segment
X25689 N25689 N25690 Segment
X25690 N25690 N25691 Segment
X25691 N25691 N25692 Segment
X25692 N25692 N25693 Segment
X25693 N25693 N25694 Segment
X25694 N25694 N25695 Segment
X25695 N25695 N25696 Segment
X25696 N25696 N25697 Segment
X25697 N25697 N25698 Segment
X25698 N25698 N25699 Segment
X25699 N25699 N25700 Segment
X25700 N25700 N25701 Segment
X25701 N25701 N25702 Segment
X25702 N25702 N25703 Segment
X25703 N25703 N25704 Segment
X25704 N25704 N25705 Segment
X25705 N25705 N25706 Segment
X25706 N25706 N25707 Segment
X25707 N25707 N25708 Segment
X25708 N25708 N25709 Segment
X25709 N25709 N25710 Segment
X25710 N25710 N25711 Segment
X25711 N25711 N25712 Segment
X25712 N25712 N25713 Segment
X25713 N25713 N25714 Segment
X25714 N25714 N25715 Segment
X25715 N25715 N25716 Segment
X25716 N25716 N25717 Segment
X25717 N25717 N25718 Segment
X25718 N25718 N25719 Segment
X25719 N25719 N25720 Segment
X25720 N25720 N25721 Segment
X25721 N25721 N25722 Segment
X25722 N25722 N25723 Segment
X25723 N25723 N25724 Segment
X25724 N25724 N25725 Segment
X25725 N25725 N25726 Segment
X25726 N25726 N25727 Segment
X25727 N25727 N25728 Segment
X25728 N25728 N25729 Segment
X25729 N25729 N25730 Segment
X25730 N25730 N25731 Segment
X25731 N25731 N25732 Segment
X25732 N25732 N25733 Segment
X25733 N25733 N25734 Segment
X25734 N25734 N25735 Segment
X25735 N25735 N25736 Segment
X25736 N25736 N25737 Segment
X25737 N25737 N25738 Segment
X25738 N25738 N25739 Segment
X25739 N25739 N25740 Segment
X25740 N25740 N25741 Segment
X25741 N25741 N25742 Segment
X25742 N25742 N25743 Segment
X25743 N25743 N25744 Segment
X25744 N25744 N25745 Segment
X25745 N25745 N25746 Segment
X25746 N25746 N25747 Segment
X25747 N25747 N25748 Segment
X25748 N25748 N25749 Segment
X25749 N25749 N25750 Segment
X25750 N25750 N25751 Segment
X25751 N25751 N25752 Segment
X25752 N25752 N25753 Segment
X25753 N25753 N25754 Segment
X25754 N25754 N25755 Segment
X25755 N25755 N25756 Segment
X25756 N25756 N25757 Segment
X25757 N25757 N25758 Segment
X25758 N25758 N25759 Segment
X25759 N25759 N25760 Segment
X25760 N25760 N25761 Segment
X25761 N25761 N25762 Segment
X25762 N25762 N25763 Segment
X25763 N25763 N25764 Segment
X25764 N25764 N25765 Segment
X25765 N25765 N25766 Segment
X25766 N25766 N25767 Segment
X25767 N25767 N25768 Segment
X25768 N25768 N25769 Segment
X25769 N25769 N25770 Segment
X25770 N25770 N25771 Segment
X25771 N25771 N25772 Segment
X25772 N25772 N25773 Segment
X25773 N25773 N25774 Segment
X25774 N25774 N25775 Segment
X25775 N25775 N25776 Segment
X25776 N25776 N25777 Segment
X25777 N25777 N25778 Segment
X25778 N25778 N25779 Segment
X25779 N25779 N25780 Segment
X25780 N25780 N25781 Segment
X25781 N25781 N25782 Segment
X25782 N25782 N25783 Segment
X25783 N25783 N25784 Segment
X25784 N25784 N25785 Segment
X25785 N25785 N25786 Segment
X25786 N25786 N25787 Segment
X25787 N25787 N25788 Segment
X25788 N25788 N25789 Segment
X25789 N25789 N25790 Segment
X25790 N25790 N25791 Segment
X25791 N25791 N25792 Segment
X25792 N25792 N25793 Segment
X25793 N25793 N25794 Segment
X25794 N25794 N25795 Segment
X25795 N25795 N25796 Segment
X25796 N25796 N25797 Segment
X25797 N25797 N25798 Segment
X25798 N25798 N25799 Segment
X25799 N25799 N25800 Segment
X25800 N25800 N25801 Segment
X25801 N25801 N25802 Segment
X25802 N25802 N25803 Segment
X25803 N25803 N25804 Segment
X25804 N25804 N25805 Segment
X25805 N25805 N25806 Segment
X25806 N25806 N25807 Segment
X25807 N25807 N25808 Segment
X25808 N25808 N25809 Segment
X25809 N25809 N25810 Segment
X25810 N25810 N25811 Segment
X25811 N25811 N25812 Segment
X25812 N25812 N25813 Segment
X25813 N25813 N25814 Segment
X25814 N25814 N25815 Segment
X25815 N25815 N25816 Segment
X25816 N25816 N25817 Segment
X25817 N25817 N25818 Segment
X25818 N25818 N25819 Segment
X25819 N25819 N25820 Segment
X25820 N25820 N25821 Segment
X25821 N25821 N25822 Segment
X25822 N25822 N25823 Segment
X25823 N25823 N25824 Segment
X25824 N25824 N25825 Segment
X25825 N25825 N25826 Segment
X25826 N25826 N25827 Segment
X25827 N25827 N25828 Segment
X25828 N25828 N25829 Segment
X25829 N25829 N25830 Segment
X25830 N25830 N25831 Segment
X25831 N25831 N25832 Segment
X25832 N25832 N25833 Segment
X25833 N25833 N25834 Segment
X25834 N25834 N25835 Segment
X25835 N25835 N25836 Segment
X25836 N25836 N25837 Segment
X25837 N25837 N25838 Segment
X25838 N25838 N25839 Segment
X25839 N25839 N25840 Segment
X25840 N25840 N25841 Segment
X25841 N25841 N25842 Segment
X25842 N25842 N25843 Segment
X25843 N25843 N25844 Segment
X25844 N25844 N25845 Segment
X25845 N25845 N25846 Segment
X25846 N25846 N25847 Segment
X25847 N25847 N25848 Segment
X25848 N25848 N25849 Segment
X25849 N25849 N25850 Segment
X25850 N25850 N25851 Segment
X25851 N25851 N25852 Segment
X25852 N25852 N25853 Segment
X25853 N25853 N25854 Segment
X25854 N25854 N25855 Segment
X25855 N25855 N25856 Segment
X25856 N25856 N25857 Segment
X25857 N25857 N25858 Segment
X25858 N25858 N25859 Segment
X25859 N25859 N25860 Segment
X25860 N25860 N25861 Segment
X25861 N25861 N25862 Segment
X25862 N25862 N25863 Segment
X25863 N25863 N25864 Segment
X25864 N25864 N25865 Segment
X25865 N25865 N25866 Segment
X25866 N25866 N25867 Segment
X25867 N25867 N25868 Segment
X25868 N25868 N25869 Segment
X25869 N25869 N25870 Segment
X25870 N25870 N25871 Segment
X25871 N25871 N25872 Segment
X25872 N25872 N25873 Segment
X25873 N25873 N25874 Segment
X25874 N25874 N25875 Segment
X25875 N25875 N25876 Segment
X25876 N25876 N25877 Segment
X25877 N25877 N25878 Segment
X25878 N25878 N25879 Segment
X25879 N25879 N25880 Segment
X25880 N25880 N25881 Segment
X25881 N25881 N25882 Segment
X25882 N25882 N25883 Segment
X25883 N25883 N25884 Segment
X25884 N25884 N25885 Segment
X25885 N25885 N25886 Segment
X25886 N25886 N25887 Segment
X25887 N25887 N25888 Segment
X25888 N25888 N25889 Segment
X25889 N25889 N25890 Segment
X25890 N25890 N25891 Segment
X25891 N25891 N25892 Segment
X25892 N25892 N25893 Segment
X25893 N25893 N25894 Segment
X25894 N25894 N25895 Segment
X25895 N25895 N25896 Segment
X25896 N25896 N25897 Segment
X25897 N25897 N25898 Segment
X25898 N25898 N25899 Segment
X25899 N25899 N25900 Segment
X25900 N25900 N25901 Segment
X25901 N25901 N25902 Segment
X25902 N25902 N25903 Segment
X25903 N25903 N25904 Segment
X25904 N25904 N25905 Segment
X25905 N25905 N25906 Segment
X25906 N25906 N25907 Segment
X25907 N25907 N25908 Segment
X25908 N25908 N25909 Segment
X25909 N25909 N25910 Segment
X25910 N25910 N25911 Segment
X25911 N25911 N25912 Segment
X25912 N25912 N25913 Segment
X25913 N25913 N25914 Segment
X25914 N25914 N25915 Segment
X25915 N25915 N25916 Segment
X25916 N25916 N25917 Segment
X25917 N25917 N25918 Segment
X25918 N25918 N25919 Segment
X25919 N25919 N25920 Segment
X25920 N25920 N25921 Segment
X25921 N25921 N25922 Segment
X25922 N25922 N25923 Segment
X25923 N25923 N25924 Segment
X25924 N25924 N25925 Segment
X25925 N25925 N25926 Segment
X25926 N25926 N25927 Segment
X25927 N25927 N25928 Segment
X25928 N25928 N25929 Segment
X25929 N25929 N25930 Segment
X25930 N25930 N25931 Segment
X25931 N25931 N25932 Segment
X25932 N25932 N25933 Segment
X25933 N25933 N25934 Segment
X25934 N25934 N25935 Segment
X25935 N25935 N25936 Segment
X25936 N25936 N25937 Segment
X25937 N25937 N25938 Segment
X25938 N25938 N25939 Segment
X25939 N25939 N25940 Segment
X25940 N25940 N25941 Segment
X25941 N25941 N25942 Segment
X25942 N25942 N25943 Segment
X25943 N25943 N25944 Segment
X25944 N25944 N25945 Segment
X25945 N25945 N25946 Segment
X25946 N25946 N25947 Segment
X25947 N25947 N25948 Segment
X25948 N25948 N25949 Segment
X25949 N25949 N25950 Segment
X25950 N25950 N25951 Segment
X25951 N25951 N25952 Segment
X25952 N25952 N25953 Segment
X25953 N25953 N25954 Segment
X25954 N25954 N25955 Segment
X25955 N25955 N25956 Segment
X25956 N25956 N25957 Segment
X25957 N25957 N25958 Segment
X25958 N25958 N25959 Segment
X25959 N25959 N25960 Segment
X25960 N25960 N25961 Segment
X25961 N25961 N25962 Segment
X25962 N25962 N25963 Segment
X25963 N25963 N25964 Segment
X25964 N25964 N25965 Segment
X25965 N25965 N25966 Segment
X25966 N25966 N25967 Segment
X25967 N25967 N25968 Segment
X25968 N25968 N25969 Segment
X25969 N25969 N25970 Segment
X25970 N25970 N25971 Segment
X25971 N25971 N25972 Segment
X25972 N25972 N25973 Segment
X25973 N25973 N25974 Segment
X25974 N25974 N25975 Segment
X25975 N25975 N25976 Segment
X25976 N25976 N25977 Segment
X25977 N25977 N25978 Segment
X25978 N25978 N25979 Segment
X25979 N25979 N25980 Segment
X25980 N25980 N25981 Segment
X25981 N25981 N25982 Segment
X25982 N25982 N25983 Segment
X25983 N25983 N25984 Segment
X25984 N25984 N25985 Segment
X25985 N25985 N25986 Segment
X25986 N25986 N25987 Segment
X25987 N25987 N25988 Segment
X25988 N25988 N25989 Segment
X25989 N25989 N25990 Segment
X25990 N25990 N25991 Segment
X25991 N25991 N25992 Segment
X25992 N25992 N25993 Segment
X25993 N25993 N25994 Segment
X25994 N25994 N25995 Segment
X25995 N25995 N25996 Segment
X25996 N25996 N25997 Segment
X25997 N25997 N25998 Segment
X25998 N25998 N25999 Segment
X25999 N25999 N26000 Segment
X26000 N26000 N26001 Segment
X26001 N26001 N26002 Segment
X26002 N26002 N26003 Segment
X26003 N26003 N26004 Segment
X26004 N26004 N26005 Segment
X26005 N26005 N26006 Segment
X26006 N26006 N26007 Segment
X26007 N26007 N26008 Segment
X26008 N26008 N26009 Segment
X26009 N26009 N26010 Segment
X26010 N26010 N26011 Segment
X26011 N26011 N26012 Segment
X26012 N26012 N26013 Segment
X26013 N26013 N26014 Segment
X26014 N26014 N26015 Segment
X26015 N26015 N26016 Segment
X26016 N26016 N26017 Segment
X26017 N26017 N26018 Segment
X26018 N26018 N26019 Segment
X26019 N26019 N26020 Segment
X26020 N26020 N26021 Segment
X26021 N26021 N26022 Segment
X26022 N26022 N26023 Segment
X26023 N26023 N26024 Segment
X26024 N26024 N26025 Segment
X26025 N26025 N26026 Segment
X26026 N26026 N26027 Segment
X26027 N26027 N26028 Segment
X26028 N26028 N26029 Segment
X26029 N26029 N26030 Segment
X26030 N26030 N26031 Segment
X26031 N26031 N26032 Segment
X26032 N26032 N26033 Segment
X26033 N26033 N26034 Segment
X26034 N26034 N26035 Segment
X26035 N26035 N26036 Segment
X26036 N26036 N26037 Segment
X26037 N26037 N26038 Segment
X26038 N26038 N26039 Segment
X26039 N26039 N26040 Segment
X26040 N26040 N26041 Segment
X26041 N26041 N26042 Segment
X26042 N26042 N26043 Segment
X26043 N26043 N26044 Segment
X26044 N26044 N26045 Segment
X26045 N26045 N26046 Segment
X26046 N26046 N26047 Segment
X26047 N26047 N26048 Segment
X26048 N26048 N26049 Segment
X26049 N26049 N26050 Segment
X26050 N26050 N26051 Segment
X26051 N26051 N26052 Segment
X26052 N26052 N26053 Segment
X26053 N26053 N26054 Segment
X26054 N26054 N26055 Segment
X26055 N26055 N26056 Segment
X26056 N26056 N26057 Segment
X26057 N26057 N26058 Segment
X26058 N26058 N26059 Segment
X26059 N26059 N26060 Segment
X26060 N26060 N26061 Segment
X26061 N26061 N26062 Segment
X26062 N26062 N26063 Segment
X26063 N26063 N26064 Segment
X26064 N26064 N26065 Segment
X26065 N26065 N26066 Segment
X26066 N26066 N26067 Segment
X26067 N26067 N26068 Segment
X26068 N26068 N26069 Segment
X26069 N26069 N26070 Segment
X26070 N26070 N26071 Segment
X26071 N26071 N26072 Segment
X26072 N26072 N26073 Segment
X26073 N26073 N26074 Segment
X26074 N26074 N26075 Segment
X26075 N26075 N26076 Segment
X26076 N26076 N26077 Segment
X26077 N26077 N26078 Segment
X26078 N26078 N26079 Segment
X26079 N26079 N26080 Segment
X26080 N26080 N26081 Segment
X26081 N26081 N26082 Segment
X26082 N26082 N26083 Segment
X26083 N26083 N26084 Segment
X26084 N26084 N26085 Segment
X26085 N26085 N26086 Segment
X26086 N26086 N26087 Segment
X26087 N26087 N26088 Segment
X26088 N26088 N26089 Segment
X26089 N26089 N26090 Segment
X26090 N26090 N26091 Segment
X26091 N26091 N26092 Segment
X26092 N26092 N26093 Segment
X26093 N26093 N26094 Segment
X26094 N26094 N26095 Segment
X26095 N26095 N26096 Segment
X26096 N26096 N26097 Segment
X26097 N26097 N26098 Segment
X26098 N26098 N26099 Segment
X26099 N26099 N26100 Segment
X26100 N26100 N26101 Segment
X26101 N26101 N26102 Segment
X26102 N26102 N26103 Segment
X26103 N26103 N26104 Segment
X26104 N26104 N26105 Segment
X26105 N26105 N26106 Segment
X26106 N26106 N26107 Segment
X26107 N26107 N26108 Segment
X26108 N26108 N26109 Segment
X26109 N26109 N26110 Segment
X26110 N26110 N26111 Segment
X26111 N26111 N26112 Segment
X26112 N26112 N26113 Segment
X26113 N26113 N26114 Segment
X26114 N26114 N26115 Segment
X26115 N26115 N26116 Segment
X26116 N26116 N26117 Segment
X26117 N26117 N26118 Segment
X26118 N26118 N26119 Segment
X26119 N26119 N26120 Segment
X26120 N26120 N26121 Segment
X26121 N26121 N26122 Segment
X26122 N26122 N26123 Segment
X26123 N26123 N26124 Segment
X26124 N26124 N26125 Segment
X26125 N26125 N26126 Segment
X26126 N26126 N26127 Segment
X26127 N26127 N26128 Segment
X26128 N26128 N26129 Segment
X26129 N26129 N26130 Segment
X26130 N26130 N26131 Segment
X26131 N26131 N26132 Segment
X26132 N26132 N26133 Segment
X26133 N26133 N26134 Segment
X26134 N26134 N26135 Segment
X26135 N26135 N26136 Segment
X26136 N26136 N26137 Segment
X26137 N26137 N26138 Segment
X26138 N26138 N26139 Segment
X26139 N26139 N26140 Segment
X26140 N26140 N26141 Segment
X26141 N26141 N26142 Segment
X26142 N26142 N26143 Segment
X26143 N26143 N26144 Segment
X26144 N26144 N26145 Segment
X26145 N26145 N26146 Segment
X26146 N26146 N26147 Segment
X26147 N26147 N26148 Segment
X26148 N26148 N26149 Segment
X26149 N26149 N26150 Segment
X26150 N26150 N26151 Segment
X26151 N26151 N26152 Segment
X26152 N26152 N26153 Segment
X26153 N26153 N26154 Segment
X26154 N26154 N26155 Segment
X26155 N26155 N26156 Segment
X26156 N26156 N26157 Segment
X26157 N26157 N26158 Segment
X26158 N26158 N26159 Segment
X26159 N26159 N26160 Segment
X26160 N26160 N26161 Segment
X26161 N26161 N26162 Segment
X26162 N26162 N26163 Segment
X26163 N26163 N26164 Segment
X26164 N26164 N26165 Segment
X26165 N26165 N26166 Segment
X26166 N26166 N26167 Segment
X26167 N26167 N26168 Segment
X26168 N26168 N26169 Segment
X26169 N26169 N26170 Segment
X26170 N26170 N26171 Segment
X26171 N26171 N26172 Segment
X26172 N26172 N26173 Segment
X26173 N26173 N26174 Segment
X26174 N26174 N26175 Segment
X26175 N26175 N26176 Segment
X26176 N26176 N26177 Segment
X26177 N26177 N26178 Segment
X26178 N26178 N26179 Segment
X26179 N26179 N26180 Segment
X26180 N26180 N26181 Segment
X26181 N26181 N26182 Segment
X26182 N26182 N26183 Segment
X26183 N26183 N26184 Segment
X26184 N26184 N26185 Segment
X26185 N26185 N26186 Segment
X26186 N26186 N26187 Segment
X26187 N26187 N26188 Segment
X26188 N26188 N26189 Segment
X26189 N26189 N26190 Segment
X26190 N26190 N26191 Segment
X26191 N26191 N26192 Segment
X26192 N26192 N26193 Segment
X26193 N26193 N26194 Segment
X26194 N26194 N26195 Segment
X26195 N26195 N26196 Segment
X26196 N26196 N26197 Segment
X26197 N26197 N26198 Segment
X26198 N26198 N26199 Segment
X26199 N26199 N26200 Segment
X26200 N26200 N26201 Segment
X26201 N26201 N26202 Segment
X26202 N26202 N26203 Segment
X26203 N26203 N26204 Segment
X26204 N26204 N26205 Segment
X26205 N26205 N26206 Segment
X26206 N26206 N26207 Segment
X26207 N26207 N26208 Segment
X26208 N26208 N26209 Segment
X26209 N26209 N26210 Segment
X26210 N26210 N26211 Segment
X26211 N26211 N26212 Segment
X26212 N26212 N26213 Segment
X26213 N26213 N26214 Segment
X26214 N26214 N26215 Segment
X26215 N26215 N26216 Segment
X26216 N26216 N26217 Segment
X26217 N26217 N26218 Segment
X26218 N26218 N26219 Segment
X26219 N26219 N26220 Segment
X26220 N26220 N26221 Segment
X26221 N26221 N26222 Segment
X26222 N26222 N26223 Segment
X26223 N26223 N26224 Segment
X26224 N26224 N26225 Segment
X26225 N26225 N26226 Segment
X26226 N26226 N26227 Segment
X26227 N26227 N26228 Segment
X26228 N26228 N26229 Segment
X26229 N26229 N26230 Segment
X26230 N26230 N26231 Segment
X26231 N26231 N26232 Segment
X26232 N26232 N26233 Segment
X26233 N26233 N26234 Segment
X26234 N26234 N26235 Segment
X26235 N26235 N26236 Segment
X26236 N26236 N26237 Segment
X26237 N26237 N26238 Segment
X26238 N26238 N26239 Segment
X26239 N26239 N26240 Segment
X26240 N26240 N26241 Segment
X26241 N26241 N26242 Segment
X26242 N26242 N26243 Segment
X26243 N26243 N26244 Segment
X26244 N26244 N26245 Segment
X26245 N26245 N26246 Segment
X26246 N26246 N26247 Segment
X26247 N26247 N26248 Segment
X26248 N26248 N26249 Segment
X26249 N26249 N26250 Segment
X26250 N26250 N26251 Segment
X26251 N26251 N26252 Segment
X26252 N26252 N26253 Segment
X26253 N26253 N26254 Segment
X26254 N26254 N26255 Segment
X26255 N26255 N26256 Segment
X26256 N26256 N26257 Segment
X26257 N26257 N26258 Segment
X26258 N26258 N26259 Segment
X26259 N26259 N26260 Segment
X26260 N26260 N26261 Segment
X26261 N26261 N26262 Segment
X26262 N26262 N26263 Segment
X26263 N26263 N26264 Segment
X26264 N26264 N26265 Segment
X26265 N26265 N26266 Segment
X26266 N26266 N26267 Segment
X26267 N26267 N26268 Segment
X26268 N26268 N26269 Segment
X26269 N26269 N26270 Segment
X26270 N26270 N26271 Segment
X26271 N26271 N26272 Segment
X26272 N26272 N26273 Segment
X26273 N26273 N26274 Segment
X26274 N26274 N26275 Segment
X26275 N26275 N26276 Segment
X26276 N26276 N26277 Segment
X26277 N26277 N26278 Segment
X26278 N26278 N26279 Segment
X26279 N26279 N26280 Segment
X26280 N26280 N26281 Segment
X26281 N26281 N26282 Segment
X26282 N26282 N26283 Segment
X26283 N26283 N26284 Segment
X26284 N26284 N26285 Segment
X26285 N26285 N26286 Segment
X26286 N26286 N26287 Segment
X26287 N26287 N26288 Segment
X26288 N26288 N26289 Segment
X26289 N26289 N26290 Segment
X26290 N26290 N26291 Segment
X26291 N26291 N26292 Segment
X26292 N26292 N26293 Segment
X26293 N26293 N26294 Segment
X26294 N26294 N26295 Segment
X26295 N26295 N26296 Segment
X26296 N26296 N26297 Segment
X26297 N26297 N26298 Segment
X26298 N26298 N26299 Segment
X26299 N26299 N26300 Segment
X26300 N26300 N26301 Segment
X26301 N26301 N26302 Segment
X26302 N26302 N26303 Segment
X26303 N26303 N26304 Segment
X26304 N26304 N26305 Segment
X26305 N26305 N26306 Segment
X26306 N26306 N26307 Segment
X26307 N26307 N26308 Segment
X26308 N26308 N26309 Segment
X26309 N26309 N26310 Segment
X26310 N26310 N26311 Segment
X26311 N26311 N26312 Segment
X26312 N26312 N26313 Segment
X26313 N26313 N26314 Segment
X26314 N26314 N26315 Segment
X26315 N26315 N26316 Segment
X26316 N26316 N26317 Segment
X26317 N26317 N26318 Segment
X26318 N26318 N26319 Segment
X26319 N26319 N26320 Segment
X26320 N26320 N26321 Segment
X26321 N26321 N26322 Segment
X26322 N26322 N26323 Segment
X26323 N26323 N26324 Segment
X26324 N26324 N26325 Segment
X26325 N26325 N26326 Segment
X26326 N26326 N26327 Segment
X26327 N26327 N26328 Segment
X26328 N26328 N26329 Segment
X26329 N26329 N26330 Segment
X26330 N26330 N26331 Segment
X26331 N26331 N26332 Segment
X26332 N26332 N26333 Segment
X26333 N26333 N26334 Segment
X26334 N26334 N26335 Segment
X26335 N26335 N26336 Segment
X26336 N26336 N26337 Segment
X26337 N26337 N26338 Segment
X26338 N26338 N26339 Segment
X26339 N26339 N26340 Segment
X26340 N26340 N26341 Segment
X26341 N26341 N26342 Segment
X26342 N26342 N26343 Segment
X26343 N26343 N26344 Segment
X26344 N26344 N26345 Segment
X26345 N26345 N26346 Segment
X26346 N26346 N26347 Segment
X26347 N26347 N26348 Segment
X26348 N26348 N26349 Segment
X26349 N26349 N26350 Segment
X26350 N26350 N26351 Segment
X26351 N26351 N26352 Segment
X26352 N26352 N26353 Segment
X26353 N26353 N26354 Segment
X26354 N26354 N26355 Segment
X26355 N26355 N26356 Segment
X26356 N26356 N26357 Segment
X26357 N26357 N26358 Segment
X26358 N26358 N26359 Segment
X26359 N26359 N26360 Segment
X26360 N26360 N26361 Segment
X26361 N26361 N26362 Segment
X26362 N26362 N26363 Segment
X26363 N26363 N26364 Segment
X26364 N26364 N26365 Segment
X26365 N26365 N26366 Segment
X26366 N26366 N26367 Segment
X26367 N26367 N26368 Segment
X26368 N26368 N26369 Segment
X26369 N26369 N26370 Segment
X26370 N26370 N26371 Segment
X26371 N26371 N26372 Segment
X26372 N26372 N26373 Segment
X26373 N26373 N26374 Segment
X26374 N26374 N26375 Segment
X26375 N26375 N26376 Segment
X26376 N26376 N26377 Segment
X26377 N26377 N26378 Segment
X26378 N26378 N26379 Segment
X26379 N26379 N26380 Segment
X26380 N26380 N26381 Segment
X26381 N26381 N26382 Segment
X26382 N26382 N26383 Segment
X26383 N26383 N26384 Segment
X26384 N26384 N26385 Segment
X26385 N26385 N26386 Segment
X26386 N26386 N26387 Segment
X26387 N26387 N26388 Segment
X26388 N26388 N26389 Segment
X26389 N26389 N26390 Segment
X26390 N26390 N26391 Segment
X26391 N26391 N26392 Segment
X26392 N26392 N26393 Segment
X26393 N26393 N26394 Segment
X26394 N26394 N26395 Segment
X26395 N26395 N26396 Segment
X26396 N26396 N26397 Segment
X26397 N26397 N26398 Segment
X26398 N26398 N26399 Segment
X26399 N26399 N26400 Segment
X26400 N26400 N26401 Segment
X26401 N26401 N26402 Segment
X26402 N26402 N26403 Segment
X26403 N26403 N26404 Segment
X26404 N26404 N26405 Segment
X26405 N26405 N26406 Segment
X26406 N26406 N26407 Segment
X26407 N26407 N26408 Segment
X26408 N26408 N26409 Segment
X26409 N26409 N26410 Segment
X26410 N26410 N26411 Segment
X26411 N26411 N26412 Segment
X26412 N26412 N26413 Segment
X26413 N26413 N26414 Segment
X26414 N26414 N26415 Segment
X26415 N26415 N26416 Segment
X26416 N26416 N26417 Segment
X26417 N26417 N26418 Segment
X26418 N26418 N26419 Segment
X26419 N26419 N26420 Segment
X26420 N26420 N26421 Segment
X26421 N26421 N26422 Segment
X26422 N26422 N26423 Segment
X26423 N26423 N26424 Segment
X26424 N26424 N26425 Segment
X26425 N26425 N26426 Segment
X26426 N26426 N26427 Segment
X26427 N26427 N26428 Segment
X26428 N26428 N26429 Segment
X26429 N26429 N26430 Segment
X26430 N26430 N26431 Segment
X26431 N26431 N26432 Segment
X26432 N26432 N26433 Segment
X26433 N26433 N26434 Segment
X26434 N26434 N26435 Segment
X26435 N26435 N26436 Segment
X26436 N26436 N26437 Segment
X26437 N26437 N26438 Segment
X26438 N26438 N26439 Segment
X26439 N26439 N26440 Segment
X26440 N26440 N26441 Segment
X26441 N26441 N26442 Segment
X26442 N26442 N26443 Segment
X26443 N26443 N26444 Segment
X26444 N26444 N26445 Segment
X26445 N26445 N26446 Segment
X26446 N26446 N26447 Segment
X26447 N26447 N26448 Segment
X26448 N26448 N26449 Segment
X26449 N26449 N26450 Segment
X26450 N26450 N26451 Segment
X26451 N26451 N26452 Segment
X26452 N26452 N26453 Segment
X26453 N26453 N26454 Segment
X26454 N26454 N26455 Segment
X26455 N26455 N26456 Segment
X26456 N26456 N26457 Segment
X26457 N26457 N26458 Segment
X26458 N26458 N26459 Segment
X26459 N26459 N26460 Segment
X26460 N26460 N26461 Segment
X26461 N26461 N26462 Segment
X26462 N26462 N26463 Segment
X26463 N26463 N26464 Segment
X26464 N26464 N26465 Segment
X26465 N26465 N26466 Segment
X26466 N26466 N26467 Segment
X26467 N26467 N26468 Segment
X26468 N26468 N26469 Segment
X26469 N26469 N26470 Segment
X26470 N26470 N26471 Segment
X26471 N26471 N26472 Segment
X26472 N26472 N26473 Segment
X26473 N26473 N26474 Segment
X26474 N26474 N26475 Segment
X26475 N26475 N26476 Segment
X26476 N26476 N26477 Segment
X26477 N26477 N26478 Segment
X26478 N26478 N26479 Segment
X26479 N26479 N26480 Segment
X26480 N26480 N26481 Segment
X26481 N26481 N26482 Segment
X26482 N26482 N26483 Segment
X26483 N26483 N26484 Segment
X26484 N26484 N26485 Segment
X26485 N26485 N26486 Segment
X26486 N26486 N26487 Segment
X26487 N26487 N26488 Segment
X26488 N26488 N26489 Segment
X26489 N26489 N26490 Segment
X26490 N26490 N26491 Segment
X26491 N26491 N26492 Segment
X26492 N26492 N26493 Segment
X26493 N26493 N26494 Segment
X26494 N26494 N26495 Segment
X26495 N26495 N26496 Segment
X26496 N26496 N26497 Segment
X26497 N26497 N26498 Segment
X26498 N26498 N26499 Segment
X26499 N26499 N26500 Segment
X26500 N26500 N26501 Segment
X26501 N26501 N26502 Segment
X26502 N26502 N26503 Segment
X26503 N26503 N26504 Segment
X26504 N26504 N26505 Segment
X26505 N26505 N26506 Segment
X26506 N26506 N26507 Segment
X26507 N26507 N26508 Segment
X26508 N26508 N26509 Segment
X26509 N26509 N26510 Segment
X26510 N26510 N26511 Segment
X26511 N26511 N26512 Segment
X26512 N26512 N26513 Segment
X26513 N26513 N26514 Segment
X26514 N26514 N26515 Segment
X26515 N26515 N26516 Segment
X26516 N26516 N26517 Segment
X26517 N26517 N26518 Segment
X26518 N26518 N26519 Segment
X26519 N26519 N26520 Segment
X26520 N26520 N26521 Segment
X26521 N26521 N26522 Segment
X26522 N26522 N26523 Segment
X26523 N26523 N26524 Segment
X26524 N26524 N26525 Segment
X26525 N26525 N26526 Segment
X26526 N26526 N26527 Segment
X26527 N26527 N26528 Segment
X26528 N26528 N26529 Segment
X26529 N26529 N26530 Segment
X26530 N26530 N26531 Segment
X26531 N26531 N26532 Segment
X26532 N26532 N26533 Segment
X26533 N26533 N26534 Segment
X26534 N26534 N26535 Segment
X26535 N26535 N26536 Segment
X26536 N26536 N26537 Segment
X26537 N26537 N26538 Segment
X26538 N26538 N26539 Segment
X26539 N26539 N26540 Segment
X26540 N26540 N26541 Segment
X26541 N26541 N26542 Segment
X26542 N26542 N26543 Segment
X26543 N26543 N26544 Segment
X26544 N26544 N26545 Segment
X26545 N26545 N26546 Segment
X26546 N26546 N26547 Segment
X26547 N26547 N26548 Segment
X26548 N26548 N26549 Segment
X26549 N26549 N26550 Segment
X26550 N26550 N26551 Segment
X26551 N26551 N26552 Segment
X26552 N26552 N26553 Segment
X26553 N26553 N26554 Segment
X26554 N26554 N26555 Segment
X26555 N26555 N26556 Segment
X26556 N26556 N26557 Segment
X26557 N26557 N26558 Segment
X26558 N26558 N26559 Segment
X26559 N26559 N26560 Segment
X26560 N26560 N26561 Segment
X26561 N26561 N26562 Segment
X26562 N26562 N26563 Segment
X26563 N26563 N26564 Segment
X26564 N26564 N26565 Segment
X26565 N26565 N26566 Segment
X26566 N26566 N26567 Segment
X26567 N26567 N26568 Segment
X26568 N26568 N26569 Segment
X26569 N26569 N26570 Segment
X26570 N26570 N26571 Segment
X26571 N26571 N26572 Segment
X26572 N26572 N26573 Segment
X26573 N26573 N26574 Segment
X26574 N26574 N26575 Segment
X26575 N26575 N26576 Segment
X26576 N26576 N26577 Segment
X26577 N26577 N26578 Segment
X26578 N26578 N26579 Segment
X26579 N26579 N26580 Segment
X26580 N26580 N26581 Segment
X26581 N26581 N26582 Segment
X26582 N26582 N26583 Segment
X26583 N26583 N26584 Segment
X26584 N26584 N26585 Segment
X26585 N26585 N26586 Segment
X26586 N26586 N26587 Segment
X26587 N26587 N26588 Segment
X26588 N26588 N26589 Segment
X26589 N26589 N26590 Segment
X26590 N26590 N26591 Segment
X26591 N26591 N26592 Segment
X26592 N26592 N26593 Segment
X26593 N26593 N26594 Segment
X26594 N26594 N26595 Segment
X26595 N26595 N26596 Segment
X26596 N26596 N26597 Segment
X26597 N26597 N26598 Segment
X26598 N26598 N26599 Segment
X26599 N26599 N26600 Segment
X26600 N26600 N26601 Segment
X26601 N26601 N26602 Segment
X26602 N26602 N26603 Segment
X26603 N26603 N26604 Segment
X26604 N26604 N26605 Segment
X26605 N26605 N26606 Segment
X26606 N26606 N26607 Segment
X26607 N26607 N26608 Segment
X26608 N26608 N26609 Segment
X26609 N26609 N26610 Segment
X26610 N26610 N26611 Segment
X26611 N26611 N26612 Segment
X26612 N26612 N26613 Segment
X26613 N26613 N26614 Segment
X26614 N26614 N26615 Segment
X26615 N26615 N26616 Segment
X26616 N26616 N26617 Segment
X26617 N26617 N26618 Segment
X26618 N26618 N26619 Segment
X26619 N26619 N26620 Segment
X26620 N26620 N26621 Segment
X26621 N26621 N26622 Segment
X26622 N26622 N26623 Segment
X26623 N26623 N26624 Segment
X26624 N26624 N26625 Segment
X26625 N26625 N26626 Segment
X26626 N26626 N26627 Segment
X26627 N26627 N26628 Segment
X26628 N26628 N26629 Segment
X26629 N26629 N26630 Segment
X26630 N26630 N26631 Segment
X26631 N26631 N26632 Segment
X26632 N26632 N26633 Segment
X26633 N26633 N26634 Segment
X26634 N26634 N26635 Segment
X26635 N26635 N26636 Segment
X26636 N26636 N26637 Segment
X26637 N26637 N26638 Segment
X26638 N26638 N26639 Segment
X26639 N26639 N26640 Segment
X26640 N26640 N26641 Segment
X26641 N26641 N26642 Segment
X26642 N26642 N26643 Segment
X26643 N26643 N26644 Segment
X26644 N26644 N26645 Segment
X26645 N26645 N26646 Segment
X26646 N26646 N26647 Segment
X26647 N26647 N26648 Segment
X26648 N26648 N26649 Segment
X26649 N26649 N26650 Segment
X26650 N26650 N26651 Segment
X26651 N26651 N26652 Segment
X26652 N26652 N26653 Segment
X26653 N26653 N26654 Segment
X26654 N26654 N26655 Segment
X26655 N26655 N26656 Segment
X26656 N26656 N26657 Segment
X26657 N26657 N26658 Segment
X26658 N26658 N26659 Segment
X26659 N26659 N26660 Segment
X26660 N26660 N26661 Segment
X26661 N26661 N26662 Segment
X26662 N26662 N26663 Segment
X26663 N26663 N26664 Segment
X26664 N26664 N26665 Segment
X26665 N26665 N26666 Segment
X26666 N26666 N26667 Segment
X26667 N26667 N26668 Segment
X26668 N26668 N26669 Segment
X26669 N26669 N26670 Segment
X26670 N26670 N26671 Segment
X26671 N26671 N26672 Segment
X26672 N26672 N26673 Segment
X26673 N26673 N26674 Segment
X26674 N26674 N26675 Segment
X26675 N26675 N26676 Segment
X26676 N26676 N26677 Segment
X26677 N26677 N26678 Segment
X26678 N26678 N26679 Segment
X26679 N26679 N26680 Segment
X26680 N26680 N26681 Segment
X26681 N26681 N26682 Segment
X26682 N26682 N26683 Segment
X26683 N26683 N26684 Segment
X26684 N26684 N26685 Segment
X26685 N26685 N26686 Segment
X26686 N26686 N26687 Segment
X26687 N26687 N26688 Segment
X26688 N26688 N26689 Segment
X26689 N26689 N26690 Segment
X26690 N26690 N26691 Segment
X26691 N26691 N26692 Segment
X26692 N26692 N26693 Segment
X26693 N26693 N26694 Segment
X26694 N26694 N26695 Segment
X26695 N26695 N26696 Segment
X26696 N26696 N26697 Segment
X26697 N26697 N26698 Segment
X26698 N26698 N26699 Segment
X26699 N26699 N26700 Segment
X26700 N26700 N26701 Segment
X26701 N26701 N26702 Segment
X26702 N26702 N26703 Segment
X26703 N26703 N26704 Segment
X26704 N26704 N26705 Segment
X26705 N26705 N26706 Segment
X26706 N26706 N26707 Segment
X26707 N26707 N26708 Segment
X26708 N26708 N26709 Segment
X26709 N26709 N26710 Segment
X26710 N26710 N26711 Segment
X26711 N26711 N26712 Segment
X26712 N26712 N26713 Segment
X26713 N26713 N26714 Segment
X26714 N26714 N26715 Segment
X26715 N26715 N26716 Segment
X26716 N26716 N26717 Segment
X26717 N26717 N26718 Segment
X26718 N26718 N26719 Segment
X26719 N26719 N26720 Segment
X26720 N26720 N26721 Segment
X26721 N26721 N26722 Segment
X26722 N26722 N26723 Segment
X26723 N26723 N26724 Segment
X26724 N26724 N26725 Segment
X26725 N26725 N26726 Segment
X26726 N26726 N26727 Segment
X26727 N26727 N26728 Segment
X26728 N26728 N26729 Segment
X26729 N26729 N26730 Segment
X26730 N26730 N26731 Segment
X26731 N26731 N26732 Segment
X26732 N26732 N26733 Segment
X26733 N26733 N26734 Segment
X26734 N26734 N26735 Segment
X26735 N26735 N26736 Segment
X26736 N26736 N26737 Segment
X26737 N26737 N26738 Segment
X26738 N26738 N26739 Segment
X26739 N26739 N26740 Segment
X26740 N26740 N26741 Segment
X26741 N26741 N26742 Segment
X26742 N26742 N26743 Segment
X26743 N26743 N26744 Segment
X26744 N26744 N26745 Segment
X26745 N26745 N26746 Segment
X26746 N26746 N26747 Segment
X26747 N26747 N26748 Segment
X26748 N26748 N26749 Segment
X26749 N26749 N26750 Segment
X26750 N26750 N26751 Segment
X26751 N26751 N26752 Segment
X26752 N26752 N26753 Segment
X26753 N26753 N26754 Segment
X26754 N26754 N26755 Segment
X26755 N26755 N26756 Segment
X26756 N26756 N26757 Segment
X26757 N26757 N26758 Segment
X26758 N26758 N26759 Segment
X26759 N26759 N26760 Segment
X26760 N26760 N26761 Segment
X26761 N26761 N26762 Segment
X26762 N26762 N26763 Segment
X26763 N26763 N26764 Segment
X26764 N26764 N26765 Segment
X26765 N26765 N26766 Segment
X26766 N26766 N26767 Segment
X26767 N26767 N26768 Segment
X26768 N26768 N26769 Segment
X26769 N26769 N26770 Segment
X26770 N26770 N26771 Segment
X26771 N26771 N26772 Segment
X26772 N26772 N26773 Segment
X26773 N26773 N26774 Segment
X26774 N26774 N26775 Segment
X26775 N26775 N26776 Segment
X26776 N26776 N26777 Segment
X26777 N26777 N26778 Segment
X26778 N26778 N26779 Segment
X26779 N26779 N26780 Segment
X26780 N26780 N26781 Segment
X26781 N26781 N26782 Segment
X26782 N26782 N26783 Segment
X26783 N26783 N26784 Segment
X26784 N26784 N26785 Segment
X26785 N26785 N26786 Segment
X26786 N26786 N26787 Segment
X26787 N26787 N26788 Segment
X26788 N26788 N26789 Segment
X26789 N26789 N26790 Segment
X26790 N26790 N26791 Segment
X26791 N26791 N26792 Segment
X26792 N26792 N26793 Segment
X26793 N26793 N26794 Segment
X26794 N26794 N26795 Segment
X26795 N26795 N26796 Segment
X26796 N26796 N26797 Segment
X26797 N26797 N26798 Segment
X26798 N26798 N26799 Segment
X26799 N26799 N26800 Segment
X26800 N26800 N26801 Segment
X26801 N26801 N26802 Segment
X26802 N26802 N26803 Segment
X26803 N26803 N26804 Segment
X26804 N26804 N26805 Segment
X26805 N26805 N26806 Segment
X26806 N26806 N26807 Segment
X26807 N26807 N26808 Segment
X26808 N26808 N26809 Segment
X26809 N26809 N26810 Segment
X26810 N26810 N26811 Segment
X26811 N26811 N26812 Segment
X26812 N26812 N26813 Segment
X26813 N26813 N26814 Segment
X26814 N26814 N26815 Segment
X26815 N26815 N26816 Segment
X26816 N26816 N26817 Segment
X26817 N26817 N26818 Segment
X26818 N26818 N26819 Segment
X26819 N26819 N26820 Segment
X26820 N26820 N26821 Segment
X26821 N26821 N26822 Segment
X26822 N26822 N26823 Segment
X26823 N26823 N26824 Segment
X26824 N26824 N26825 Segment
X26825 N26825 N26826 Segment
X26826 N26826 N26827 Segment
X26827 N26827 N26828 Segment
X26828 N26828 N26829 Segment
X26829 N26829 N26830 Segment
X26830 N26830 N26831 Segment
X26831 N26831 N26832 Segment
X26832 N26832 N26833 Segment
X26833 N26833 N26834 Segment
X26834 N26834 N26835 Segment
X26835 N26835 N26836 Segment
X26836 N26836 N26837 Segment
X26837 N26837 N26838 Segment
X26838 N26838 N26839 Segment
X26839 N26839 N26840 Segment
X26840 N26840 N26841 Segment
X26841 N26841 N26842 Segment
X26842 N26842 N26843 Segment
X26843 N26843 N26844 Segment
X26844 N26844 N26845 Segment
X26845 N26845 N26846 Segment
X26846 N26846 N26847 Segment
X26847 N26847 N26848 Segment
X26848 N26848 N26849 Segment
X26849 N26849 N26850 Segment
X26850 N26850 N26851 Segment
X26851 N26851 N26852 Segment
X26852 N26852 N26853 Segment
X26853 N26853 N26854 Segment
X26854 N26854 N26855 Segment
X26855 N26855 N26856 Segment
X26856 N26856 N26857 Segment
X26857 N26857 N26858 Segment
X26858 N26858 N26859 Segment
X26859 N26859 N26860 Segment
X26860 N26860 N26861 Segment
X26861 N26861 N26862 Segment
X26862 N26862 N26863 Segment
X26863 N26863 N26864 Segment
X26864 N26864 N26865 Segment
X26865 N26865 N26866 Segment
X26866 N26866 N26867 Segment
X26867 N26867 N26868 Segment
X26868 N26868 N26869 Segment
X26869 N26869 N26870 Segment
X26870 N26870 N26871 Segment
X26871 N26871 N26872 Segment
X26872 N26872 N26873 Segment
X26873 N26873 N26874 Segment
X26874 N26874 N26875 Segment
X26875 N26875 N26876 Segment
X26876 N26876 N26877 Segment
X26877 N26877 N26878 Segment
X26878 N26878 N26879 Segment
X26879 N26879 N26880 Segment
X26880 N26880 N26881 Segment
X26881 N26881 N26882 Segment
X26882 N26882 N26883 Segment
X26883 N26883 N26884 Segment
X26884 N26884 N26885 Segment
X26885 N26885 N26886 Segment
X26886 N26886 N26887 Segment
X26887 N26887 N26888 Segment
X26888 N26888 N26889 Segment
X26889 N26889 N26890 Segment
X26890 N26890 N26891 Segment
X26891 N26891 N26892 Segment
X26892 N26892 N26893 Segment
X26893 N26893 N26894 Segment
X26894 N26894 N26895 Segment
X26895 N26895 N26896 Segment
X26896 N26896 N26897 Segment
X26897 N26897 N26898 Segment
X26898 N26898 N26899 Segment
X26899 N26899 N26900 Segment
X26900 N26900 N26901 Segment
X26901 N26901 N26902 Segment
X26902 N26902 N26903 Segment
X26903 N26903 N26904 Segment
X26904 N26904 N26905 Segment
X26905 N26905 N26906 Segment
X26906 N26906 N26907 Segment
X26907 N26907 N26908 Segment
X26908 N26908 N26909 Segment
X26909 N26909 N26910 Segment
X26910 N26910 N26911 Segment
X26911 N26911 N26912 Segment
X26912 N26912 N26913 Segment
X26913 N26913 N26914 Segment
X26914 N26914 N26915 Segment
X26915 N26915 N26916 Segment
X26916 N26916 N26917 Segment
X26917 N26917 N26918 Segment
X26918 N26918 N26919 Segment
X26919 N26919 N26920 Segment
X26920 N26920 N26921 Segment
X26921 N26921 N26922 Segment
X26922 N26922 N26923 Segment
X26923 N26923 N26924 Segment
X26924 N26924 N26925 Segment
X26925 N26925 N26926 Segment
X26926 N26926 N26927 Segment
X26927 N26927 N26928 Segment
X26928 N26928 N26929 Segment
X26929 N26929 N26930 Segment
X26930 N26930 N26931 Segment
X26931 N26931 N26932 Segment
X26932 N26932 N26933 Segment
X26933 N26933 N26934 Segment
X26934 N26934 N26935 Segment
X26935 N26935 N26936 Segment
X26936 N26936 N26937 Segment
X26937 N26937 N26938 Segment
X26938 N26938 N26939 Segment
X26939 N26939 N26940 Segment
X26940 N26940 N26941 Segment
X26941 N26941 N26942 Segment
X26942 N26942 N26943 Segment
X26943 N26943 N26944 Segment
X26944 N26944 N26945 Segment
X26945 N26945 N26946 Segment
X26946 N26946 N26947 Segment
X26947 N26947 N26948 Segment
X26948 N26948 N26949 Segment
X26949 N26949 N26950 Segment
X26950 N26950 N26951 Segment
X26951 N26951 N26952 Segment
X26952 N26952 N26953 Segment
X26953 N26953 N26954 Segment
X26954 N26954 N26955 Segment
X26955 N26955 N26956 Segment
X26956 N26956 N26957 Segment
X26957 N26957 N26958 Segment
X26958 N26958 N26959 Segment
X26959 N26959 N26960 Segment
X26960 N26960 N26961 Segment
X26961 N26961 N26962 Segment
X26962 N26962 N26963 Segment
X26963 N26963 N26964 Segment
X26964 N26964 N26965 Segment
X26965 N26965 N26966 Segment
X26966 N26966 N26967 Segment
X26967 N26967 N26968 Segment
X26968 N26968 N26969 Segment
X26969 N26969 N26970 Segment
X26970 N26970 N26971 Segment
X26971 N26971 N26972 Segment
X26972 N26972 N26973 Segment
X26973 N26973 N26974 Segment
X26974 N26974 N26975 Segment
X26975 N26975 N26976 Segment
X26976 N26976 N26977 Segment
X26977 N26977 N26978 Segment
X26978 N26978 N26979 Segment
X26979 N26979 N26980 Segment
X26980 N26980 N26981 Segment
X26981 N26981 N26982 Segment
X26982 N26982 N26983 Segment
X26983 N26983 N26984 Segment
X26984 N26984 N26985 Segment
X26985 N26985 N26986 Segment
X26986 N26986 N26987 Segment
X26987 N26987 N26988 Segment
X26988 N26988 N26989 Segment
X26989 N26989 N26990 Segment
X26990 N26990 N26991 Segment
X26991 N26991 N26992 Segment
X26992 N26992 N26993 Segment
X26993 N26993 N26994 Segment
X26994 N26994 N26995 Segment
X26995 N26995 N26996 Segment
X26996 N26996 N26997 Segment
X26997 N26997 N26998 Segment
X26998 N26998 N26999 Segment
X26999 N26999 N27000 Segment
X27000 N27000 N27001 Segment
X27001 N27001 N27002 Segment
X27002 N27002 N27003 Segment
X27003 N27003 N27004 Segment
X27004 N27004 N27005 Segment
X27005 N27005 N27006 Segment
X27006 N27006 N27007 Segment
X27007 N27007 N27008 Segment
X27008 N27008 N27009 Segment
X27009 N27009 N27010 Segment
X27010 N27010 N27011 Segment
X27011 N27011 N27012 Segment
X27012 N27012 N27013 Segment
X27013 N27013 N27014 Segment
X27014 N27014 N27015 Segment
X27015 N27015 N27016 Segment
X27016 N27016 N27017 Segment
X27017 N27017 N27018 Segment
X27018 N27018 N27019 Segment
X27019 N27019 N27020 Segment
X27020 N27020 N27021 Segment
X27021 N27021 N27022 Segment
X27022 N27022 N27023 Segment
X27023 N27023 N27024 Segment
X27024 N27024 N27025 Segment
X27025 N27025 N27026 Segment
X27026 N27026 N27027 Segment
X27027 N27027 N27028 Segment
X27028 N27028 N27029 Segment
X27029 N27029 N27030 Segment
X27030 N27030 N27031 Segment
X27031 N27031 N27032 Segment
X27032 N27032 N27033 Segment
X27033 N27033 N27034 Segment
X27034 N27034 N27035 Segment
X27035 N27035 N27036 Segment
X27036 N27036 N27037 Segment
X27037 N27037 N27038 Segment
X27038 N27038 N27039 Segment
X27039 N27039 N27040 Segment
X27040 N27040 N27041 Segment
X27041 N27041 N27042 Segment
X27042 N27042 N27043 Segment
X27043 N27043 N27044 Segment
X27044 N27044 N27045 Segment
X27045 N27045 N27046 Segment
X27046 N27046 N27047 Segment
X27047 N27047 N27048 Segment
X27048 N27048 N27049 Segment
X27049 N27049 N27050 Segment
X27050 N27050 N27051 Segment
X27051 N27051 N27052 Segment
X27052 N27052 N27053 Segment
X27053 N27053 N27054 Segment
X27054 N27054 N27055 Segment
X27055 N27055 N27056 Segment
X27056 N27056 N27057 Segment
X27057 N27057 N27058 Segment
X27058 N27058 N27059 Segment
X27059 N27059 N27060 Segment
X27060 N27060 N27061 Segment
X27061 N27061 N27062 Segment
X27062 N27062 N27063 Segment
X27063 N27063 N27064 Segment
X27064 N27064 N27065 Segment
X27065 N27065 N27066 Segment
X27066 N27066 N27067 Segment
X27067 N27067 N27068 Segment
X27068 N27068 N27069 Segment
X27069 N27069 N27070 Segment
X27070 N27070 N27071 Segment
X27071 N27071 N27072 Segment
X27072 N27072 N27073 Segment
X27073 N27073 N27074 Segment
X27074 N27074 N27075 Segment
X27075 N27075 N27076 Segment
X27076 N27076 N27077 Segment
X27077 N27077 N27078 Segment
X27078 N27078 N27079 Segment
X27079 N27079 N27080 Segment
X27080 N27080 N27081 Segment
X27081 N27081 N27082 Segment
X27082 N27082 N27083 Segment
X27083 N27083 N27084 Segment
X27084 N27084 N27085 Segment
X27085 N27085 N27086 Segment
X27086 N27086 N27087 Segment
X27087 N27087 N27088 Segment
X27088 N27088 N27089 Segment
X27089 N27089 N27090 Segment
X27090 N27090 N27091 Segment
X27091 N27091 N27092 Segment
X27092 N27092 N27093 Segment
X27093 N27093 N27094 Segment
X27094 N27094 N27095 Segment
X27095 N27095 N27096 Segment
X27096 N27096 N27097 Segment
X27097 N27097 N27098 Segment
X27098 N27098 N27099 Segment
X27099 N27099 N27100 Segment
X27100 N27100 N27101 Segment
X27101 N27101 N27102 Segment
X27102 N27102 N27103 Segment
X27103 N27103 N27104 Segment
X27104 N27104 N27105 Segment
X27105 N27105 N27106 Segment
X27106 N27106 N27107 Segment
X27107 N27107 N27108 Segment
X27108 N27108 N27109 Segment
X27109 N27109 N27110 Segment
X27110 N27110 N27111 Segment
X27111 N27111 N27112 Segment
X27112 N27112 N27113 Segment
X27113 N27113 N27114 Segment
X27114 N27114 N27115 Segment
X27115 N27115 N27116 Segment
X27116 N27116 N27117 Segment
X27117 N27117 N27118 Segment
X27118 N27118 N27119 Segment
X27119 N27119 N27120 Segment
X27120 N27120 N27121 Segment
X27121 N27121 N27122 Segment
X27122 N27122 N27123 Segment
X27123 N27123 N27124 Segment
X27124 N27124 N27125 Segment
X27125 N27125 N27126 Segment
X27126 N27126 N27127 Segment
X27127 N27127 N27128 Segment
X27128 N27128 N27129 Segment
X27129 N27129 N27130 Segment
X27130 N27130 N27131 Segment
X27131 N27131 N27132 Segment
X27132 N27132 N27133 Segment
X27133 N27133 N27134 Segment
X27134 N27134 N27135 Segment
X27135 N27135 N27136 Segment
X27136 N27136 N27137 Segment
X27137 N27137 N27138 Segment
X27138 N27138 N27139 Segment
X27139 N27139 N27140 Segment
X27140 N27140 N27141 Segment
X27141 N27141 N27142 Segment
X27142 N27142 N27143 Segment
X27143 N27143 N27144 Segment
X27144 N27144 N27145 Segment
X27145 N27145 N27146 Segment
X27146 N27146 N27147 Segment
X27147 N27147 N27148 Segment
X27148 N27148 N27149 Segment
X27149 N27149 N27150 Segment
X27150 N27150 N27151 Segment
X27151 N27151 N27152 Segment
X27152 N27152 N27153 Segment
X27153 N27153 N27154 Segment
X27154 N27154 N27155 Segment
X27155 N27155 N27156 Segment
X27156 N27156 N27157 Segment
X27157 N27157 N27158 Segment
X27158 N27158 N27159 Segment
X27159 N27159 N27160 Segment
X27160 N27160 N27161 Segment
X27161 N27161 N27162 Segment
X27162 N27162 N27163 Segment
X27163 N27163 N27164 Segment
X27164 N27164 N27165 Segment
X27165 N27165 N27166 Segment
X27166 N27166 N27167 Segment
X27167 N27167 N27168 Segment
X27168 N27168 N27169 Segment
X27169 N27169 N27170 Segment
X27170 N27170 N27171 Segment
X27171 N27171 N27172 Segment
X27172 N27172 N27173 Segment
X27173 N27173 N27174 Segment
X27174 N27174 N27175 Segment
X27175 N27175 N27176 Segment
X27176 N27176 N27177 Segment
X27177 N27177 N27178 Segment
X27178 N27178 N27179 Segment
X27179 N27179 N27180 Segment
X27180 N27180 N27181 Segment
X27181 N27181 N27182 Segment
X27182 N27182 N27183 Segment
X27183 N27183 N27184 Segment
X27184 N27184 N27185 Segment
X27185 N27185 N27186 Segment
X27186 N27186 N27187 Segment
X27187 N27187 N27188 Segment
X27188 N27188 N27189 Segment
X27189 N27189 N27190 Segment
X27190 N27190 N27191 Segment
X27191 N27191 N27192 Segment
X27192 N27192 N27193 Segment
X27193 N27193 N27194 Segment
X27194 N27194 N27195 Segment
X27195 N27195 N27196 Segment
X27196 N27196 N27197 Segment
X27197 N27197 N27198 Segment
X27198 N27198 N27199 Segment
X27199 N27199 N27200 Segment
X27200 N27200 N27201 Segment
X27201 N27201 N27202 Segment
X27202 N27202 N27203 Segment
X27203 N27203 N27204 Segment
X27204 N27204 N27205 Segment
X27205 N27205 N27206 Segment
X27206 N27206 N27207 Segment
X27207 N27207 N27208 Segment
X27208 N27208 N27209 Segment
X27209 N27209 N27210 Segment
X27210 N27210 N27211 Segment
X27211 N27211 N27212 Segment
X27212 N27212 N27213 Segment
X27213 N27213 N27214 Segment
X27214 N27214 N27215 Segment
X27215 N27215 N27216 Segment
X27216 N27216 N27217 Segment
X27217 N27217 N27218 Segment
X27218 N27218 N27219 Segment
X27219 N27219 N27220 Segment
X27220 N27220 N27221 Segment
X27221 N27221 N27222 Segment
X27222 N27222 N27223 Segment
X27223 N27223 N27224 Segment
X27224 N27224 N27225 Segment
X27225 N27225 N27226 Segment
X27226 N27226 N27227 Segment
X27227 N27227 N27228 Segment
X27228 N27228 N27229 Segment
X27229 N27229 N27230 Segment
X27230 N27230 N27231 Segment
X27231 N27231 N27232 Segment
X27232 N27232 N27233 Segment
X27233 N27233 N27234 Segment
X27234 N27234 N27235 Segment
X27235 N27235 N27236 Segment
X27236 N27236 N27237 Segment
X27237 N27237 N27238 Segment
X27238 N27238 N27239 Segment
X27239 N27239 N27240 Segment
X27240 N27240 N27241 Segment
X27241 N27241 N27242 Segment
X27242 N27242 N27243 Segment
X27243 N27243 N27244 Segment
X27244 N27244 N27245 Segment
X27245 N27245 N27246 Segment
X27246 N27246 N27247 Segment
X27247 N27247 N27248 Segment
X27248 N27248 N27249 Segment
X27249 N27249 N27250 Segment
X27250 N27250 N27251 Segment
X27251 N27251 N27252 Segment
X27252 N27252 N27253 Segment
X27253 N27253 N27254 Segment
X27254 N27254 N27255 Segment
X27255 N27255 N27256 Segment
X27256 N27256 N27257 Segment
X27257 N27257 N27258 Segment
X27258 N27258 N27259 Segment
X27259 N27259 N27260 Segment
X27260 N27260 N27261 Segment
X27261 N27261 N27262 Segment
X27262 N27262 N27263 Segment
X27263 N27263 N27264 Segment
X27264 N27264 N27265 Segment
X27265 N27265 N27266 Segment
X27266 N27266 N27267 Segment
X27267 N27267 N27268 Segment
X27268 N27268 N27269 Segment
X27269 N27269 N27270 Segment
X27270 N27270 N27271 Segment
X27271 N27271 N27272 Segment
X27272 N27272 N27273 Segment
X27273 N27273 N27274 Segment
X27274 N27274 N27275 Segment
X27275 N27275 N27276 Segment
X27276 N27276 N27277 Segment
X27277 N27277 N27278 Segment
X27278 N27278 N27279 Segment
X27279 N27279 N27280 Segment
X27280 N27280 N27281 Segment
X27281 N27281 N27282 Segment
X27282 N27282 N27283 Segment
X27283 N27283 N27284 Segment
X27284 N27284 N27285 Segment
X27285 N27285 N27286 Segment
X27286 N27286 N27287 Segment
X27287 N27287 N27288 Segment
X27288 N27288 N27289 Segment
X27289 N27289 N27290 Segment
X27290 N27290 N27291 Segment
X27291 N27291 N27292 Segment
X27292 N27292 N27293 Segment
X27293 N27293 N27294 Segment
X27294 N27294 N27295 Segment
X27295 N27295 N27296 Segment
X27296 N27296 N27297 Segment
X27297 N27297 N27298 Segment
X27298 N27298 N27299 Segment
X27299 N27299 N27300 Segment
X27300 N27300 N27301 Segment
X27301 N27301 N27302 Segment
X27302 N27302 N27303 Segment
X27303 N27303 N27304 Segment
X27304 N27304 N27305 Segment
X27305 N27305 N27306 Segment
X27306 N27306 N27307 Segment
X27307 N27307 N27308 Segment
X27308 N27308 N27309 Segment
X27309 N27309 N27310 Segment
X27310 N27310 N27311 Segment
X27311 N27311 N27312 Segment
X27312 N27312 N27313 Segment
X27313 N27313 N27314 Segment
X27314 N27314 N27315 Segment
X27315 N27315 N27316 Segment
X27316 N27316 N27317 Segment
X27317 N27317 N27318 Segment
X27318 N27318 N27319 Segment
X27319 N27319 N27320 Segment
X27320 N27320 N27321 Segment
X27321 N27321 N27322 Segment
X27322 N27322 N27323 Segment
X27323 N27323 N27324 Segment
X27324 N27324 N27325 Segment
X27325 N27325 N27326 Segment
X27326 N27326 N27327 Segment
X27327 N27327 N27328 Segment
X27328 N27328 N27329 Segment
X27329 N27329 N27330 Segment
X27330 N27330 N27331 Segment
X27331 N27331 N27332 Segment
X27332 N27332 N27333 Segment
X27333 N27333 N27334 Segment
X27334 N27334 N27335 Segment
X27335 N27335 N27336 Segment
X27336 N27336 N27337 Segment
X27337 N27337 N27338 Segment
X27338 N27338 N27339 Segment
X27339 N27339 N27340 Segment
X27340 N27340 N27341 Segment
X27341 N27341 N27342 Segment
X27342 N27342 N27343 Segment
X27343 N27343 N27344 Segment
X27344 N27344 N27345 Segment
X27345 N27345 N27346 Segment
X27346 N27346 N27347 Segment
X27347 N27347 N27348 Segment
X27348 N27348 N27349 Segment
X27349 N27349 N27350 Segment
X27350 N27350 N27351 Segment
X27351 N27351 N27352 Segment
X27352 N27352 N27353 Segment
X27353 N27353 N27354 Segment
X27354 N27354 N27355 Segment
X27355 N27355 N27356 Segment
X27356 N27356 N27357 Segment
X27357 N27357 N27358 Segment
X27358 N27358 N27359 Segment
X27359 N27359 N27360 Segment
X27360 N27360 N27361 Segment
X27361 N27361 N27362 Segment
X27362 N27362 N27363 Segment
X27363 N27363 N27364 Segment
X27364 N27364 N27365 Segment
X27365 N27365 N27366 Segment
X27366 N27366 N27367 Segment
X27367 N27367 N27368 Segment
X27368 N27368 N27369 Segment
X27369 N27369 N27370 Segment
X27370 N27370 N27371 Segment
X27371 N27371 N27372 Segment
X27372 N27372 N27373 Segment
X27373 N27373 N27374 Segment
X27374 N27374 N27375 Segment
X27375 N27375 N27376 Segment
X27376 N27376 N27377 Segment
X27377 N27377 N27378 Segment
X27378 N27378 N27379 Segment
X27379 N27379 N27380 Segment
X27380 N27380 N27381 Segment
X27381 N27381 N27382 Segment
X27382 N27382 N27383 Segment
X27383 N27383 N27384 Segment
X27384 N27384 N27385 Segment
X27385 N27385 N27386 Segment
X27386 N27386 N27387 Segment
X27387 N27387 N27388 Segment
X27388 N27388 N27389 Segment
X27389 N27389 N27390 Segment
X27390 N27390 N27391 Segment
X27391 N27391 N27392 Segment
X27392 N27392 N27393 Segment
X27393 N27393 N27394 Segment
X27394 N27394 N27395 Segment
X27395 N27395 N27396 Segment
X27396 N27396 N27397 Segment
X27397 N27397 N27398 Segment
X27398 N27398 N27399 Segment
X27399 N27399 N27400 Segment
X27400 N27400 N27401 Segment
X27401 N27401 N27402 Segment
X27402 N27402 N27403 Segment
X27403 N27403 N27404 Segment
X27404 N27404 N27405 Segment
X27405 N27405 N27406 Segment
X27406 N27406 N27407 Segment
X27407 N27407 N27408 Segment
X27408 N27408 N27409 Segment
X27409 N27409 N27410 Segment
X27410 N27410 N27411 Segment
X27411 N27411 N27412 Segment
X27412 N27412 N27413 Segment
X27413 N27413 N27414 Segment
X27414 N27414 N27415 Segment
X27415 N27415 N27416 Segment
X27416 N27416 N27417 Segment
X27417 N27417 N27418 Segment
X27418 N27418 N27419 Segment
X27419 N27419 N27420 Segment
X27420 N27420 N27421 Segment
X27421 N27421 N27422 Segment
X27422 N27422 N27423 Segment
X27423 N27423 N27424 Segment
X27424 N27424 N27425 Segment
X27425 N27425 N27426 Segment
X27426 N27426 N27427 Segment
X27427 N27427 N27428 Segment
X27428 N27428 N27429 Segment
X27429 N27429 N27430 Segment
X27430 N27430 N27431 Segment
X27431 N27431 N27432 Segment
X27432 N27432 N27433 Segment
X27433 N27433 N27434 Segment
X27434 N27434 N27435 Segment
X27435 N27435 N27436 Segment
X27436 N27436 N27437 Segment
X27437 N27437 N27438 Segment
X27438 N27438 N27439 Segment
X27439 N27439 N27440 Segment
X27440 N27440 N27441 Segment
X27441 N27441 N27442 Segment
X27442 N27442 N27443 Segment
X27443 N27443 N27444 Segment
X27444 N27444 N27445 Segment
X27445 N27445 N27446 Segment
X27446 N27446 N27447 Segment
X27447 N27447 N27448 Segment
X27448 N27448 N27449 Segment
X27449 N27449 N27450 Segment
X27450 N27450 N27451 Segment
X27451 N27451 N27452 Segment
X27452 N27452 N27453 Segment
X27453 N27453 N27454 Segment
X27454 N27454 N27455 Segment
X27455 N27455 N27456 Segment
X27456 N27456 N27457 Segment
X27457 N27457 N27458 Segment
X27458 N27458 N27459 Segment
X27459 N27459 N27460 Segment
X27460 N27460 N27461 Segment
X27461 N27461 N27462 Segment
X27462 N27462 N27463 Segment
X27463 N27463 N27464 Segment
X27464 N27464 N27465 Segment
X27465 N27465 N27466 Segment
X27466 N27466 N27467 Segment
X27467 N27467 N27468 Segment
X27468 N27468 N27469 Segment
X27469 N27469 N27470 Segment
X27470 N27470 N27471 Segment
X27471 N27471 N27472 Segment
X27472 N27472 N27473 Segment
X27473 N27473 N27474 Segment
X27474 N27474 N27475 Segment
X27475 N27475 N27476 Segment
X27476 N27476 N27477 Segment
X27477 N27477 N27478 Segment
X27478 N27478 N27479 Segment
X27479 N27479 N27480 Segment
X27480 N27480 N27481 Segment
X27481 N27481 N27482 Segment
X27482 N27482 N27483 Segment
X27483 N27483 N27484 Segment
X27484 N27484 N27485 Segment
X27485 N27485 N27486 Segment
X27486 N27486 N27487 Segment
X27487 N27487 N27488 Segment
X27488 N27488 N27489 Segment
X27489 N27489 N27490 Segment
X27490 N27490 N27491 Segment
X27491 N27491 N27492 Segment
X27492 N27492 N27493 Segment
X27493 N27493 N27494 Segment
X27494 N27494 N27495 Segment
X27495 N27495 N27496 Segment
X27496 N27496 N27497 Segment
X27497 N27497 N27498 Segment
X27498 N27498 N27499 Segment
X27499 N27499 N27500 Segment
X27500 N27500 N27501 Segment
X27501 N27501 N27502 Segment
X27502 N27502 N27503 Segment
X27503 N27503 N27504 Segment
X27504 N27504 N27505 Segment
X27505 N27505 N27506 Segment
X27506 N27506 N27507 Segment
X27507 N27507 N27508 Segment
X27508 N27508 N27509 Segment
X27509 N27509 N27510 Segment
X27510 N27510 N27511 Segment
X27511 N27511 N27512 Segment
X27512 N27512 N27513 Segment
X27513 N27513 N27514 Segment
X27514 N27514 N27515 Segment
X27515 N27515 N27516 Segment
X27516 N27516 N27517 Segment
X27517 N27517 N27518 Segment
X27518 N27518 N27519 Segment
X27519 N27519 N27520 Segment
X27520 N27520 N27521 Segment
X27521 N27521 N27522 Segment
X27522 N27522 N27523 Segment
X27523 N27523 N27524 Segment
X27524 N27524 N27525 Segment
X27525 N27525 N27526 Segment
X27526 N27526 N27527 Segment
X27527 N27527 N27528 Segment
X27528 N27528 N27529 Segment
X27529 N27529 N27530 Segment
X27530 N27530 N27531 Segment
X27531 N27531 N27532 Segment
X27532 N27532 N27533 Segment
X27533 N27533 N27534 Segment
X27534 N27534 N27535 Segment
X27535 N27535 N27536 Segment
X27536 N27536 N27537 Segment
X27537 N27537 N27538 Segment
X27538 N27538 N27539 Segment
X27539 N27539 N27540 Segment
X27540 N27540 N27541 Segment
X27541 N27541 N27542 Segment
X27542 N27542 N27543 Segment
X27543 N27543 N27544 Segment
X27544 N27544 N27545 Segment
X27545 N27545 N27546 Segment
X27546 N27546 N27547 Segment
X27547 N27547 N27548 Segment
X27548 N27548 N27549 Segment
X27549 N27549 N27550 Segment
X27550 N27550 N27551 Segment
X27551 N27551 N27552 Segment
X27552 N27552 N27553 Segment
X27553 N27553 N27554 Segment
X27554 N27554 N27555 Segment
X27555 N27555 N27556 Segment
X27556 N27556 N27557 Segment
X27557 N27557 N27558 Segment
X27558 N27558 N27559 Segment
X27559 N27559 N27560 Segment
X27560 N27560 N27561 Segment
X27561 N27561 N27562 Segment
X27562 N27562 N27563 Segment
X27563 N27563 N27564 Segment
X27564 N27564 N27565 Segment
X27565 N27565 N27566 Segment
X27566 N27566 N27567 Segment
X27567 N27567 N27568 Segment
X27568 N27568 N27569 Segment
X27569 N27569 N27570 Segment
X27570 N27570 N27571 Segment
X27571 N27571 N27572 Segment
X27572 N27572 N27573 Segment
X27573 N27573 N27574 Segment
X27574 N27574 N27575 Segment
X27575 N27575 N27576 Segment
X27576 N27576 N27577 Segment
X27577 N27577 N27578 Segment
X27578 N27578 N27579 Segment
X27579 N27579 N27580 Segment
X27580 N27580 N27581 Segment
X27581 N27581 N27582 Segment
X27582 N27582 N27583 Segment
X27583 N27583 N27584 Segment
X27584 N27584 N27585 Segment
X27585 N27585 N27586 Segment
X27586 N27586 N27587 Segment
X27587 N27587 N27588 Segment
X27588 N27588 N27589 Segment
X27589 N27589 N27590 Segment
X27590 N27590 N27591 Segment
X27591 N27591 N27592 Segment
X27592 N27592 N27593 Segment
X27593 N27593 N27594 Segment
X27594 N27594 N27595 Segment
X27595 N27595 N27596 Segment
X27596 N27596 N27597 Segment
X27597 N27597 N27598 Segment
X27598 N27598 N27599 Segment
X27599 N27599 N27600 Segment
X27600 N27600 N27601 Segment
X27601 N27601 N27602 Segment
X27602 N27602 N27603 Segment
X27603 N27603 N27604 Segment
X27604 N27604 N27605 Segment
X27605 N27605 N27606 Segment
X27606 N27606 N27607 Segment
X27607 N27607 N27608 Segment
X27608 N27608 N27609 Segment
X27609 N27609 N27610 Segment
X27610 N27610 N27611 Segment
X27611 N27611 N27612 Segment
X27612 N27612 N27613 Segment
X27613 N27613 N27614 Segment
X27614 N27614 N27615 Segment
X27615 N27615 N27616 Segment
X27616 N27616 N27617 Segment
X27617 N27617 N27618 Segment
X27618 N27618 N27619 Segment
X27619 N27619 N27620 Segment
X27620 N27620 N27621 Segment
X27621 N27621 N27622 Segment
X27622 N27622 N27623 Segment
X27623 N27623 N27624 Segment
X27624 N27624 N27625 Segment
X27625 N27625 N27626 Segment
X27626 N27626 N27627 Segment
X27627 N27627 N27628 Segment
X27628 N27628 N27629 Segment
X27629 N27629 N27630 Segment
X27630 N27630 N27631 Segment
X27631 N27631 N27632 Segment
X27632 N27632 N27633 Segment
X27633 N27633 N27634 Segment
X27634 N27634 N27635 Segment
X27635 N27635 N27636 Segment
X27636 N27636 N27637 Segment
X27637 N27637 N27638 Segment
X27638 N27638 N27639 Segment
X27639 N27639 N27640 Segment
X27640 N27640 N27641 Segment
X27641 N27641 N27642 Segment
X27642 N27642 N27643 Segment
X27643 N27643 N27644 Segment
X27644 N27644 N27645 Segment
X27645 N27645 N27646 Segment
X27646 N27646 N27647 Segment
X27647 N27647 N27648 Segment
X27648 N27648 N27649 Segment
X27649 N27649 N27650 Segment
X27650 N27650 N27651 Segment
X27651 N27651 N27652 Segment
X27652 N27652 N27653 Segment
X27653 N27653 N27654 Segment
X27654 N27654 N27655 Segment
X27655 N27655 N27656 Segment
X27656 N27656 N27657 Segment
X27657 N27657 N27658 Segment
X27658 N27658 N27659 Segment
X27659 N27659 N27660 Segment
X27660 N27660 N27661 Segment
X27661 N27661 N27662 Segment
X27662 N27662 N27663 Segment
X27663 N27663 N27664 Segment
X27664 N27664 N27665 Segment
X27665 N27665 N27666 Segment
X27666 N27666 N27667 Segment
X27667 N27667 N27668 Segment
X27668 N27668 N27669 Segment
X27669 N27669 N27670 Segment
X27670 N27670 N27671 Segment
X27671 N27671 N27672 Segment
X27672 N27672 N27673 Segment
X27673 N27673 N27674 Segment
X27674 N27674 N27675 Segment
X27675 N27675 N27676 Segment
X27676 N27676 N27677 Segment
X27677 N27677 N27678 Segment
X27678 N27678 N27679 Segment
X27679 N27679 N27680 Segment
X27680 N27680 N27681 Segment
X27681 N27681 N27682 Segment
X27682 N27682 N27683 Segment
X27683 N27683 N27684 Segment
X27684 N27684 N27685 Segment
X27685 N27685 N27686 Segment
X27686 N27686 N27687 Segment
X27687 N27687 N27688 Segment
X27688 N27688 N27689 Segment
X27689 N27689 N27690 Segment
X27690 N27690 N27691 Segment
X27691 N27691 N27692 Segment
X27692 N27692 N27693 Segment
X27693 N27693 N27694 Segment
X27694 N27694 N27695 Segment
X27695 N27695 N27696 Segment
X27696 N27696 N27697 Segment
X27697 N27697 N27698 Segment
X27698 N27698 N27699 Segment
X27699 N27699 N27700 Segment
X27700 N27700 N27701 Segment
X27701 N27701 N27702 Segment
X27702 N27702 N27703 Segment
X27703 N27703 N27704 Segment
X27704 N27704 N27705 Segment
X27705 N27705 N27706 Segment
X27706 N27706 N27707 Segment
X27707 N27707 N27708 Segment
X27708 N27708 N27709 Segment
X27709 N27709 N27710 Segment
X27710 N27710 N27711 Segment
X27711 N27711 N27712 Segment
X27712 N27712 N27713 Segment
X27713 N27713 N27714 Segment
X27714 N27714 N27715 Segment
X27715 N27715 N27716 Segment
X27716 N27716 N27717 Segment
X27717 N27717 N27718 Segment
X27718 N27718 N27719 Segment
X27719 N27719 N27720 Segment
X27720 N27720 N27721 Segment
X27721 N27721 N27722 Segment
X27722 N27722 N27723 Segment
X27723 N27723 N27724 Segment
X27724 N27724 N27725 Segment
X27725 N27725 N27726 Segment
X27726 N27726 N27727 Segment
X27727 N27727 N27728 Segment
X27728 N27728 N27729 Segment
X27729 N27729 N27730 Segment
X27730 N27730 N27731 Segment
X27731 N27731 N27732 Segment
X27732 N27732 N27733 Segment
X27733 N27733 N27734 Segment
X27734 N27734 N27735 Segment
X27735 N27735 N27736 Segment
X27736 N27736 N27737 Segment
X27737 N27737 N27738 Segment
X27738 N27738 N27739 Segment
X27739 N27739 N27740 Segment
X27740 N27740 N27741 Segment
X27741 N27741 N27742 Segment
X27742 N27742 N27743 Segment
X27743 N27743 N27744 Segment
X27744 N27744 N27745 Segment
X27745 N27745 N27746 Segment
X27746 N27746 N27747 Segment
X27747 N27747 N27748 Segment
X27748 N27748 N27749 Segment
X27749 N27749 N27750 Segment
X27750 N27750 N27751 Segment
X27751 N27751 N27752 Segment
X27752 N27752 N27753 Segment
X27753 N27753 N27754 Segment
X27754 N27754 N27755 Segment
X27755 N27755 N27756 Segment
X27756 N27756 N27757 Segment
X27757 N27757 N27758 Segment
X27758 N27758 N27759 Segment
X27759 N27759 N27760 Segment
X27760 N27760 N27761 Segment
X27761 N27761 N27762 Segment
X27762 N27762 N27763 Segment
X27763 N27763 N27764 Segment
X27764 N27764 N27765 Segment
X27765 N27765 N27766 Segment
X27766 N27766 N27767 Segment
X27767 N27767 N27768 Segment
X27768 N27768 N27769 Segment
X27769 N27769 N27770 Segment
X27770 N27770 N27771 Segment
X27771 N27771 N27772 Segment
X27772 N27772 N27773 Segment
X27773 N27773 N27774 Segment
X27774 N27774 N27775 Segment
X27775 N27775 N27776 Segment
X27776 N27776 N27777 Segment
X27777 N27777 N27778 Segment
X27778 N27778 N27779 Segment
X27779 N27779 N27780 Segment
X27780 N27780 N27781 Segment
X27781 N27781 N27782 Segment
X27782 N27782 N27783 Segment
X27783 N27783 N27784 Segment
X27784 N27784 N27785 Segment
X27785 N27785 N27786 Segment
X27786 N27786 N27787 Segment
X27787 N27787 N27788 Segment
X27788 N27788 N27789 Segment
X27789 N27789 N27790 Segment
X27790 N27790 N27791 Segment
X27791 N27791 N27792 Segment
X27792 N27792 N27793 Segment
X27793 N27793 N27794 Segment
X27794 N27794 N27795 Segment
X27795 N27795 N27796 Segment
X27796 N27796 N27797 Segment
X27797 N27797 N27798 Segment
X27798 N27798 N27799 Segment
X27799 N27799 N27800 Segment
X27800 N27800 N27801 Segment
X27801 N27801 N27802 Segment
X27802 N27802 N27803 Segment
X27803 N27803 N27804 Segment
X27804 N27804 N27805 Segment
X27805 N27805 N27806 Segment
X27806 N27806 N27807 Segment
X27807 N27807 N27808 Segment
X27808 N27808 N27809 Segment
X27809 N27809 N27810 Segment
X27810 N27810 N27811 Segment
X27811 N27811 N27812 Segment
X27812 N27812 N27813 Segment
X27813 N27813 N27814 Segment
X27814 N27814 N27815 Segment
X27815 N27815 N27816 Segment
X27816 N27816 N27817 Segment
X27817 N27817 N27818 Segment
X27818 N27818 N27819 Segment
X27819 N27819 N27820 Segment
X27820 N27820 N27821 Segment
X27821 N27821 N27822 Segment
X27822 N27822 N27823 Segment
X27823 N27823 N27824 Segment
X27824 N27824 N27825 Segment
X27825 N27825 N27826 Segment
X27826 N27826 N27827 Segment
X27827 N27827 N27828 Segment
X27828 N27828 N27829 Segment
X27829 N27829 N27830 Segment
X27830 N27830 N27831 Segment
X27831 N27831 N27832 Segment
X27832 N27832 N27833 Segment
X27833 N27833 N27834 Segment
X27834 N27834 N27835 Segment
X27835 N27835 N27836 Segment
X27836 N27836 N27837 Segment
X27837 N27837 N27838 Segment
X27838 N27838 N27839 Segment
X27839 N27839 N27840 Segment
X27840 N27840 N27841 Segment
X27841 N27841 N27842 Segment
X27842 N27842 N27843 Segment
X27843 N27843 N27844 Segment
X27844 N27844 N27845 Segment
X27845 N27845 N27846 Segment
X27846 N27846 N27847 Segment
X27847 N27847 N27848 Segment
X27848 N27848 N27849 Segment
X27849 N27849 N27850 Segment
X27850 N27850 N27851 Segment
X27851 N27851 N27852 Segment
X27852 N27852 N27853 Segment
X27853 N27853 N27854 Segment
X27854 N27854 N27855 Segment
X27855 N27855 N27856 Segment
X27856 N27856 N27857 Segment
X27857 N27857 N27858 Segment
X27858 N27858 N27859 Segment
X27859 N27859 N27860 Segment
X27860 N27860 N27861 Segment
X27861 N27861 N27862 Segment
X27862 N27862 N27863 Segment
X27863 N27863 N27864 Segment
X27864 N27864 N27865 Segment
X27865 N27865 N27866 Segment
X27866 N27866 N27867 Segment
X27867 N27867 N27868 Segment
X27868 N27868 N27869 Segment
X27869 N27869 N27870 Segment
X27870 N27870 N27871 Segment
X27871 N27871 N27872 Segment
X27872 N27872 N27873 Segment
X27873 N27873 N27874 Segment
X27874 N27874 N27875 Segment
X27875 N27875 N27876 Segment
X27876 N27876 N27877 Segment
X27877 N27877 N27878 Segment
X27878 N27878 N27879 Segment
X27879 N27879 N27880 Segment
X27880 N27880 N27881 Segment
X27881 N27881 N27882 Segment
X27882 N27882 N27883 Segment
X27883 N27883 N27884 Segment
X27884 N27884 N27885 Segment
X27885 N27885 N27886 Segment
X27886 N27886 N27887 Segment
X27887 N27887 N27888 Segment
X27888 N27888 N27889 Segment
X27889 N27889 N27890 Segment
X27890 N27890 N27891 Segment
X27891 N27891 N27892 Segment
X27892 N27892 N27893 Segment
X27893 N27893 N27894 Segment
X27894 N27894 N27895 Segment
X27895 N27895 N27896 Segment
X27896 N27896 N27897 Segment
X27897 N27897 N27898 Segment
X27898 N27898 N27899 Segment
X27899 N27899 N27900 Segment
X27900 N27900 N27901 Segment
X27901 N27901 N27902 Segment
X27902 N27902 N27903 Segment
X27903 N27903 N27904 Segment
X27904 N27904 N27905 Segment
X27905 N27905 N27906 Segment
X27906 N27906 N27907 Segment
X27907 N27907 N27908 Segment
X27908 N27908 N27909 Segment
X27909 N27909 N27910 Segment
X27910 N27910 N27911 Segment
X27911 N27911 N27912 Segment
X27912 N27912 N27913 Segment
X27913 N27913 N27914 Segment
X27914 N27914 N27915 Segment
X27915 N27915 N27916 Segment
X27916 N27916 N27917 Segment
X27917 N27917 N27918 Segment
X27918 N27918 N27919 Segment
X27919 N27919 N27920 Segment
X27920 N27920 N27921 Segment
X27921 N27921 N27922 Segment
X27922 N27922 N27923 Segment
X27923 N27923 N27924 Segment
X27924 N27924 N27925 Segment
X27925 N27925 N27926 Segment
X27926 N27926 N27927 Segment
X27927 N27927 N27928 Segment
X27928 N27928 N27929 Segment
X27929 N27929 N27930 Segment
X27930 N27930 N27931 Segment
X27931 N27931 N27932 Segment
X27932 N27932 N27933 Segment
X27933 N27933 N27934 Segment
X27934 N27934 N27935 Segment
X27935 N27935 N27936 Segment
X27936 N27936 N27937 Segment
X27937 N27937 N27938 Segment
X27938 N27938 N27939 Segment
X27939 N27939 N27940 Segment
X27940 N27940 N27941 Segment
X27941 N27941 N27942 Segment
X27942 N27942 N27943 Segment
X27943 N27943 N27944 Segment
X27944 N27944 N27945 Segment
X27945 N27945 N27946 Segment
X27946 N27946 N27947 Segment
X27947 N27947 N27948 Segment
X27948 N27948 N27949 Segment
X27949 N27949 N27950 Segment
X27950 N27950 N27951 Segment
X27951 N27951 N27952 Segment
X27952 N27952 N27953 Segment
X27953 N27953 N27954 Segment
X27954 N27954 N27955 Segment
X27955 N27955 N27956 Segment
X27956 N27956 N27957 Segment
X27957 N27957 N27958 Segment
X27958 N27958 N27959 Segment
X27959 N27959 N27960 Segment
X27960 N27960 N27961 Segment
X27961 N27961 N27962 Segment
X27962 N27962 N27963 Segment
X27963 N27963 N27964 Segment
X27964 N27964 N27965 Segment
X27965 N27965 N27966 Segment
X27966 N27966 N27967 Segment
X27967 N27967 N27968 Segment
X27968 N27968 N27969 Segment
X27969 N27969 N27970 Segment
X27970 N27970 N27971 Segment
X27971 N27971 N27972 Segment
X27972 N27972 N27973 Segment
X27973 N27973 N27974 Segment
X27974 N27974 N27975 Segment
X27975 N27975 N27976 Segment
X27976 N27976 N27977 Segment
X27977 N27977 N27978 Segment
X27978 N27978 N27979 Segment
X27979 N27979 N27980 Segment
X27980 N27980 N27981 Segment
X27981 N27981 N27982 Segment
X27982 N27982 N27983 Segment
X27983 N27983 N27984 Segment
X27984 N27984 N27985 Segment
X27985 N27985 N27986 Segment
X27986 N27986 N27987 Segment
X27987 N27987 N27988 Segment
X27988 N27988 N27989 Segment
X27989 N27989 N27990 Segment
X27990 N27990 N27991 Segment
X27991 N27991 N27992 Segment
X27992 N27992 N27993 Segment
X27993 N27993 N27994 Segment
X27994 N27994 N27995 Segment
X27995 N27995 N27996 Segment
X27996 N27996 N27997 Segment
X27997 N27997 N27998 Segment
X27998 N27998 N27999 Segment
X27999 N27999 N28000 Segment
X28000 N28000 N28001 Segment
X28001 N28001 N28002 Segment
X28002 N28002 N28003 Segment
X28003 N28003 N28004 Segment
X28004 N28004 N28005 Segment
X28005 N28005 N28006 Segment
X28006 N28006 N28007 Segment
X28007 N28007 N28008 Segment
X28008 N28008 N28009 Segment
X28009 N28009 N28010 Segment
X28010 N28010 N28011 Segment
X28011 N28011 N28012 Segment
X28012 N28012 N28013 Segment
X28013 N28013 N28014 Segment
X28014 N28014 N28015 Segment
X28015 N28015 N28016 Segment
X28016 N28016 N28017 Segment
X28017 N28017 N28018 Segment
X28018 N28018 N28019 Segment
X28019 N28019 N28020 Segment
X28020 N28020 N28021 Segment
X28021 N28021 N28022 Segment
X28022 N28022 N28023 Segment
X28023 N28023 N28024 Segment
X28024 N28024 N28025 Segment
X28025 N28025 N28026 Segment
X28026 N28026 N28027 Segment
X28027 N28027 N28028 Segment
X28028 N28028 N28029 Segment
X28029 N28029 N28030 Segment
X28030 N28030 N28031 Segment
X28031 N28031 N28032 Segment
X28032 N28032 N28033 Segment
X28033 N28033 N28034 Segment
X28034 N28034 N28035 Segment
X28035 N28035 N28036 Segment
X28036 N28036 N28037 Segment
X28037 N28037 N28038 Segment
X28038 N28038 N28039 Segment
X28039 N28039 N28040 Segment
X28040 N28040 N28041 Segment
X28041 N28041 N28042 Segment
X28042 N28042 N28043 Segment
X28043 N28043 N28044 Segment
X28044 N28044 N28045 Segment
X28045 N28045 N28046 Segment
X28046 N28046 N28047 Segment
X28047 N28047 N28048 Segment
X28048 N28048 N28049 Segment
X28049 N28049 N28050 Segment
X28050 N28050 N28051 Segment
X28051 N28051 N28052 Segment
X28052 N28052 N28053 Segment
X28053 N28053 N28054 Segment
X28054 N28054 N28055 Segment
X28055 N28055 N28056 Segment
X28056 N28056 N28057 Segment
X28057 N28057 N28058 Segment
X28058 N28058 N28059 Segment
X28059 N28059 N28060 Segment
X28060 N28060 N28061 Segment
X28061 N28061 N28062 Segment
X28062 N28062 N28063 Segment
X28063 N28063 N28064 Segment
X28064 N28064 N28065 Segment
X28065 N28065 N28066 Segment
X28066 N28066 N28067 Segment
X28067 N28067 N28068 Segment
X28068 N28068 N28069 Segment
X28069 N28069 N28070 Segment
X28070 N28070 N28071 Segment
X28071 N28071 N28072 Segment
X28072 N28072 N28073 Segment
X28073 N28073 N28074 Segment
X28074 N28074 N28075 Segment
X28075 N28075 N28076 Segment
X28076 N28076 N28077 Segment
X28077 N28077 N28078 Segment
X28078 N28078 N28079 Segment
X28079 N28079 N28080 Segment
X28080 N28080 N28081 Segment
X28081 N28081 N28082 Segment
X28082 N28082 N28083 Segment
X28083 N28083 N28084 Segment
X28084 N28084 N28085 Segment
X28085 N28085 N28086 Segment
X28086 N28086 N28087 Segment
X28087 N28087 N28088 Segment
X28088 N28088 N28089 Segment
X28089 N28089 N28090 Segment
X28090 N28090 N28091 Segment
X28091 N28091 N28092 Segment
X28092 N28092 N28093 Segment
X28093 N28093 N28094 Segment
X28094 N28094 N28095 Segment
X28095 N28095 N28096 Segment
X28096 N28096 N28097 Segment
X28097 N28097 N28098 Segment
X28098 N28098 N28099 Segment
X28099 N28099 N28100 Segment
X28100 N28100 N28101 Segment
X28101 N28101 N28102 Segment
X28102 N28102 N28103 Segment
X28103 N28103 N28104 Segment
X28104 N28104 N28105 Segment
X28105 N28105 N28106 Segment
X28106 N28106 N28107 Segment
X28107 N28107 N28108 Segment
X28108 N28108 N28109 Segment
X28109 N28109 N28110 Segment
X28110 N28110 N28111 Segment
X28111 N28111 N28112 Segment
X28112 N28112 N28113 Segment
X28113 N28113 N28114 Segment
X28114 N28114 N28115 Segment
X28115 N28115 N28116 Segment
X28116 N28116 N28117 Segment
X28117 N28117 N28118 Segment
X28118 N28118 N28119 Segment
X28119 N28119 N28120 Segment
X28120 N28120 N28121 Segment
X28121 N28121 N28122 Segment
X28122 N28122 N28123 Segment
X28123 N28123 N28124 Segment
X28124 N28124 N28125 Segment
X28125 N28125 N28126 Segment
X28126 N28126 N28127 Segment
X28127 N28127 N28128 Segment
X28128 N28128 N28129 Segment
X28129 N28129 N28130 Segment
X28130 N28130 N28131 Segment
X28131 N28131 N28132 Segment
X28132 N28132 N28133 Segment
X28133 N28133 N28134 Segment
X28134 N28134 N28135 Segment
X28135 N28135 N28136 Segment
X28136 N28136 N28137 Segment
X28137 N28137 N28138 Segment
X28138 N28138 N28139 Segment
X28139 N28139 N28140 Segment
X28140 N28140 N28141 Segment
X28141 N28141 N28142 Segment
X28142 N28142 N28143 Segment
X28143 N28143 N28144 Segment
X28144 N28144 N28145 Segment
X28145 N28145 N28146 Segment
X28146 N28146 N28147 Segment
X28147 N28147 N28148 Segment
X28148 N28148 N28149 Segment
X28149 N28149 N28150 Segment
X28150 N28150 N28151 Segment
X28151 N28151 N28152 Segment
X28152 N28152 N28153 Segment
X28153 N28153 N28154 Segment
X28154 N28154 N28155 Segment
X28155 N28155 N28156 Segment
X28156 N28156 N28157 Segment
X28157 N28157 N28158 Segment
X28158 N28158 N28159 Segment
X28159 N28159 N28160 Segment
X28160 N28160 N28161 Segment
X28161 N28161 N28162 Segment
X28162 N28162 N28163 Segment
X28163 N28163 N28164 Segment
X28164 N28164 N28165 Segment
X28165 N28165 N28166 Segment
X28166 N28166 N28167 Segment
X28167 N28167 N28168 Segment
X28168 N28168 N28169 Segment
X28169 N28169 N28170 Segment
X28170 N28170 N28171 Segment
X28171 N28171 N28172 Segment
X28172 N28172 N28173 Segment
X28173 N28173 N28174 Segment
X28174 N28174 N28175 Segment
X28175 N28175 N28176 Segment
X28176 N28176 N28177 Segment
X28177 N28177 N28178 Segment
X28178 N28178 N28179 Segment
X28179 N28179 N28180 Segment
X28180 N28180 N28181 Segment
X28181 N28181 N28182 Segment
X28182 N28182 N28183 Segment
X28183 N28183 N28184 Segment
X28184 N28184 N28185 Segment
X28185 N28185 N28186 Segment
X28186 N28186 N28187 Segment
X28187 N28187 N28188 Segment
X28188 N28188 N28189 Segment
X28189 N28189 N28190 Segment
X28190 N28190 N28191 Segment
X28191 N28191 N28192 Segment
X28192 N28192 N28193 Segment
X28193 N28193 N28194 Segment
X28194 N28194 N28195 Segment
X28195 N28195 N28196 Segment
X28196 N28196 N28197 Segment
X28197 N28197 N28198 Segment
X28198 N28198 N28199 Segment
X28199 N28199 N28200 Segment
X28200 N28200 N28201 Segment
X28201 N28201 N28202 Segment
X28202 N28202 N28203 Segment
X28203 N28203 N28204 Segment
X28204 N28204 N28205 Segment
X28205 N28205 N28206 Segment
X28206 N28206 N28207 Segment
X28207 N28207 N28208 Segment
X28208 N28208 N28209 Segment
X28209 N28209 N28210 Segment
X28210 N28210 N28211 Segment
X28211 N28211 N28212 Segment
X28212 N28212 N28213 Segment
X28213 N28213 N28214 Segment
X28214 N28214 N28215 Segment
X28215 N28215 N28216 Segment
X28216 N28216 N28217 Segment
X28217 N28217 N28218 Segment
X28218 N28218 N28219 Segment
X28219 N28219 N28220 Segment
X28220 N28220 N28221 Segment
X28221 N28221 N28222 Segment
X28222 N28222 N28223 Segment
X28223 N28223 N28224 Segment
X28224 N28224 N28225 Segment
X28225 N28225 N28226 Segment
X28226 N28226 N28227 Segment
X28227 N28227 N28228 Segment
X28228 N28228 N28229 Segment
X28229 N28229 N28230 Segment
X28230 N28230 N28231 Segment
X28231 N28231 N28232 Segment
X28232 N28232 N28233 Segment
X28233 N28233 N28234 Segment
X28234 N28234 N28235 Segment
X28235 N28235 N28236 Segment
X28236 N28236 N28237 Segment
X28237 N28237 N28238 Segment
X28238 N28238 N28239 Segment
X28239 N28239 N28240 Segment
X28240 N28240 N28241 Segment
X28241 N28241 N28242 Segment
X28242 N28242 N28243 Segment
X28243 N28243 N28244 Segment
X28244 N28244 N28245 Segment
X28245 N28245 N28246 Segment
X28246 N28246 N28247 Segment
X28247 N28247 N28248 Segment
X28248 N28248 N28249 Segment
X28249 N28249 N28250 Segment
X28250 N28250 N28251 Segment
X28251 N28251 N28252 Segment
X28252 N28252 N28253 Segment
X28253 N28253 N28254 Segment
X28254 N28254 N28255 Segment
X28255 N28255 N28256 Segment
X28256 N28256 N28257 Segment
X28257 N28257 N28258 Segment
X28258 N28258 N28259 Segment
X28259 N28259 N28260 Segment
X28260 N28260 N28261 Segment
X28261 N28261 N28262 Segment
X28262 N28262 N28263 Segment
X28263 N28263 N28264 Segment
X28264 N28264 N28265 Segment
X28265 N28265 N28266 Segment
X28266 N28266 N28267 Segment
X28267 N28267 N28268 Segment
X28268 N28268 N28269 Segment
X28269 N28269 N28270 Segment
X28270 N28270 N28271 Segment
X28271 N28271 N28272 Segment
X28272 N28272 N28273 Segment
X28273 N28273 N28274 Segment
X28274 N28274 N28275 Segment
X28275 N28275 N28276 Segment
X28276 N28276 N28277 Segment
X28277 N28277 N28278 Segment
X28278 N28278 N28279 Segment
X28279 N28279 N28280 Segment
X28280 N28280 N28281 Segment
X28281 N28281 N28282 Segment
X28282 N28282 N28283 Segment
X28283 N28283 N28284 Segment
X28284 N28284 N28285 Segment
X28285 N28285 N28286 Segment
X28286 N28286 N28287 Segment
X28287 N28287 N28288 Segment
X28288 N28288 N28289 Segment
X28289 N28289 N28290 Segment
X28290 N28290 N28291 Segment
X28291 N28291 N28292 Segment
X28292 N28292 N28293 Segment
X28293 N28293 N28294 Segment
X28294 N28294 N28295 Segment
X28295 N28295 N28296 Segment
X28296 N28296 N28297 Segment
X28297 N28297 N28298 Segment
X28298 N28298 N28299 Segment
X28299 N28299 N28300 Segment
X28300 N28300 N28301 Segment
X28301 N28301 N28302 Segment
X28302 N28302 N28303 Segment
X28303 N28303 N28304 Segment
X28304 N28304 N28305 Segment
X28305 N28305 N28306 Segment
X28306 N28306 N28307 Segment
X28307 N28307 N28308 Segment
X28308 N28308 N28309 Segment
X28309 N28309 N28310 Segment
X28310 N28310 N28311 Segment
X28311 N28311 N28312 Segment
X28312 N28312 N28313 Segment
X28313 N28313 N28314 Segment
X28314 N28314 N28315 Segment
X28315 N28315 N28316 Segment
X28316 N28316 N28317 Segment
X28317 N28317 N28318 Segment
X28318 N28318 N28319 Segment
X28319 N28319 N28320 Segment
X28320 N28320 N28321 Segment
X28321 N28321 N28322 Segment
X28322 N28322 N28323 Segment
X28323 N28323 N28324 Segment
X28324 N28324 N28325 Segment
X28325 N28325 N28326 Segment
X28326 N28326 N28327 Segment
X28327 N28327 N28328 Segment
X28328 N28328 N28329 Segment
X28329 N28329 N28330 Segment
X28330 N28330 N28331 Segment
X28331 N28331 N28332 Segment
X28332 N28332 N28333 Segment
X28333 N28333 N28334 Segment
X28334 N28334 N28335 Segment
X28335 N28335 N28336 Segment
X28336 N28336 N28337 Segment
X28337 N28337 N28338 Segment
X28338 N28338 N28339 Segment
X28339 N28339 N28340 Segment
X28340 N28340 N28341 Segment
X28341 N28341 N28342 Segment
X28342 N28342 N28343 Segment
X28343 N28343 N28344 Segment
X28344 N28344 N28345 Segment
X28345 N28345 N28346 Segment
X28346 N28346 N28347 Segment
X28347 N28347 N28348 Segment
X28348 N28348 N28349 Segment
X28349 N28349 N28350 Segment
X28350 N28350 N28351 Segment
X28351 N28351 N28352 Segment
X28352 N28352 N28353 Segment
X28353 N28353 N28354 Segment
X28354 N28354 N28355 Segment
X28355 N28355 N28356 Segment
X28356 N28356 N28357 Segment
X28357 N28357 N28358 Segment
X28358 N28358 N28359 Segment
X28359 N28359 N28360 Segment
X28360 N28360 N28361 Segment
X28361 N28361 N28362 Segment
X28362 N28362 N28363 Segment
X28363 N28363 N28364 Segment
X28364 N28364 N28365 Segment
X28365 N28365 N28366 Segment
X28366 N28366 N28367 Segment
X28367 N28367 N28368 Segment
X28368 N28368 N28369 Segment
X28369 N28369 N28370 Segment
X28370 N28370 N28371 Segment
X28371 N28371 N28372 Segment
X28372 N28372 N28373 Segment
X28373 N28373 N28374 Segment
X28374 N28374 N28375 Segment
X28375 N28375 N28376 Segment
X28376 N28376 N28377 Segment
X28377 N28377 N28378 Segment
X28378 N28378 N28379 Segment
X28379 N28379 N28380 Segment
X28380 N28380 N28381 Segment
X28381 N28381 N28382 Segment
X28382 N28382 N28383 Segment
X28383 N28383 N28384 Segment
X28384 N28384 N28385 Segment
X28385 N28385 N28386 Segment
X28386 N28386 N28387 Segment
X28387 N28387 N28388 Segment
X28388 N28388 N28389 Segment
X28389 N28389 N28390 Segment
X28390 N28390 N28391 Segment
X28391 N28391 N28392 Segment
X28392 N28392 N28393 Segment
X28393 N28393 N28394 Segment
X28394 N28394 N28395 Segment
X28395 N28395 N28396 Segment
X28396 N28396 N28397 Segment
X28397 N28397 N28398 Segment
X28398 N28398 N28399 Segment
X28399 N28399 N28400 Segment
X28400 N28400 N28401 Segment
X28401 N28401 N28402 Segment
X28402 N28402 N28403 Segment
X28403 N28403 N28404 Segment
X28404 N28404 N28405 Segment
X28405 N28405 N28406 Segment
X28406 N28406 N28407 Segment
X28407 N28407 N28408 Segment
X28408 N28408 N28409 Segment
X28409 N28409 N28410 Segment
X28410 N28410 N28411 Segment
X28411 N28411 N28412 Segment
X28412 N28412 N28413 Segment
X28413 N28413 N28414 Segment
X28414 N28414 N28415 Segment
X28415 N28415 N28416 Segment
X28416 N28416 N28417 Segment
X28417 N28417 N28418 Segment
X28418 N28418 N28419 Segment
X28419 N28419 N28420 Segment
X28420 N28420 N28421 Segment
X28421 N28421 N28422 Segment
X28422 N28422 N28423 Segment
X28423 N28423 N28424 Segment
X28424 N28424 N28425 Segment
X28425 N28425 N28426 Segment
X28426 N28426 N28427 Segment
X28427 N28427 N28428 Segment
X28428 N28428 N28429 Segment
X28429 N28429 N28430 Segment
X28430 N28430 N28431 Segment
X28431 N28431 N28432 Segment
X28432 N28432 N28433 Segment
X28433 N28433 N28434 Segment
X28434 N28434 N28435 Segment
X28435 N28435 N28436 Segment
X28436 N28436 N28437 Segment
X28437 N28437 N28438 Segment
X28438 N28438 N28439 Segment
X28439 N28439 N28440 Segment
X28440 N28440 N28441 Segment
X28441 N28441 N28442 Segment
X28442 N28442 N28443 Segment
X28443 N28443 N28444 Segment
X28444 N28444 N28445 Segment
X28445 N28445 N28446 Segment
X28446 N28446 N28447 Segment
X28447 N28447 N28448 Segment
X28448 N28448 N28449 Segment
X28449 N28449 N28450 Segment
X28450 N28450 N28451 Segment
X28451 N28451 N28452 Segment
X28452 N28452 N28453 Segment
X28453 N28453 N28454 Segment
X28454 N28454 N28455 Segment
X28455 N28455 N28456 Segment
X28456 N28456 N28457 Segment
X28457 N28457 N28458 Segment
X28458 N28458 N28459 Segment
X28459 N28459 N28460 Segment
X28460 N28460 N28461 Segment
X28461 N28461 N28462 Segment
X28462 N28462 N28463 Segment
X28463 N28463 N28464 Segment
X28464 N28464 N28465 Segment
X28465 N28465 N28466 Segment
X28466 N28466 N28467 Segment
X28467 N28467 N28468 Segment
X28468 N28468 N28469 Segment
X28469 N28469 N28470 Segment
X28470 N28470 N28471 Segment
X28471 N28471 N28472 Segment
X28472 N28472 N28473 Segment
X28473 N28473 N28474 Segment
X28474 N28474 N28475 Segment
X28475 N28475 N28476 Segment
X28476 N28476 N28477 Segment
X28477 N28477 N28478 Segment
X28478 N28478 N28479 Segment
X28479 N28479 N28480 Segment
X28480 N28480 N28481 Segment
X28481 N28481 N28482 Segment
X28482 N28482 N28483 Segment
X28483 N28483 N28484 Segment
X28484 N28484 N28485 Segment
X28485 N28485 N28486 Segment
X28486 N28486 N28487 Segment
X28487 N28487 N28488 Segment
X28488 N28488 N28489 Segment
X28489 N28489 N28490 Segment
X28490 N28490 N28491 Segment
X28491 N28491 N28492 Segment
X28492 N28492 N28493 Segment
X28493 N28493 N28494 Segment
X28494 N28494 N28495 Segment
X28495 N28495 N28496 Segment
X28496 N28496 N28497 Segment
X28497 N28497 N28498 Segment
X28498 N28498 N28499 Segment
X28499 N28499 N28500 Segment
X28500 N28500 N28501 Segment
X28501 N28501 N28502 Segment
X28502 N28502 N28503 Segment
X28503 N28503 N28504 Segment
X28504 N28504 N28505 Segment
X28505 N28505 N28506 Segment
X28506 N28506 N28507 Segment
X28507 N28507 N28508 Segment
X28508 N28508 N28509 Segment
X28509 N28509 N28510 Segment
X28510 N28510 N28511 Segment
X28511 N28511 N28512 Segment
X28512 N28512 N28513 Segment
X28513 N28513 N28514 Segment
X28514 N28514 N28515 Segment
X28515 N28515 N28516 Segment
X28516 N28516 N28517 Segment
X28517 N28517 N28518 Segment
X28518 N28518 N28519 Segment
X28519 N28519 N28520 Segment
X28520 N28520 N28521 Segment
X28521 N28521 N28522 Segment
X28522 N28522 N28523 Segment
X28523 N28523 N28524 Segment
X28524 N28524 N28525 Segment
X28525 N28525 N28526 Segment
X28526 N28526 N28527 Segment
X28527 N28527 N28528 Segment
X28528 N28528 N28529 Segment
X28529 N28529 N28530 Segment
X28530 N28530 N28531 Segment
X28531 N28531 N28532 Segment
X28532 N28532 N28533 Segment
X28533 N28533 N28534 Segment
X28534 N28534 N28535 Segment
X28535 N28535 N28536 Segment
X28536 N28536 N28537 Segment
X28537 N28537 N28538 Segment
X28538 N28538 N28539 Segment
X28539 N28539 N28540 Segment
X28540 N28540 N28541 Segment
X28541 N28541 N28542 Segment
X28542 N28542 N28543 Segment
X28543 N28543 N28544 Segment
X28544 N28544 N28545 Segment
X28545 N28545 N28546 Segment
X28546 N28546 N28547 Segment
X28547 N28547 N28548 Segment
X28548 N28548 N28549 Segment
X28549 N28549 N28550 Segment
X28550 N28550 N28551 Segment
X28551 N28551 N28552 Segment
X28552 N28552 N28553 Segment
X28553 N28553 N28554 Segment
X28554 N28554 N28555 Segment
X28555 N28555 N28556 Segment
X28556 N28556 N28557 Segment
X28557 N28557 N28558 Segment
X28558 N28558 N28559 Segment
X28559 N28559 N28560 Segment
X28560 N28560 N28561 Segment
X28561 N28561 N28562 Segment
X28562 N28562 N28563 Segment
X28563 N28563 N28564 Segment
X28564 N28564 N28565 Segment
X28565 N28565 N28566 Segment
X28566 N28566 N28567 Segment
X28567 N28567 N28568 Segment
X28568 N28568 N28569 Segment
X28569 N28569 N28570 Segment
X28570 N28570 N28571 Segment
X28571 N28571 N28572 Segment
X28572 N28572 N28573 Segment
X28573 N28573 N28574 Segment
X28574 N28574 N28575 Segment
X28575 N28575 N28576 Segment
X28576 N28576 N28577 Segment
X28577 N28577 N28578 Segment
X28578 N28578 N28579 Segment
X28579 N28579 N28580 Segment
X28580 N28580 N28581 Segment
X28581 N28581 N28582 Segment
X28582 N28582 N28583 Segment
X28583 N28583 N28584 Segment
X28584 N28584 N28585 Segment
X28585 N28585 N28586 Segment
X28586 N28586 N28587 Segment
X28587 N28587 N28588 Segment
X28588 N28588 N28589 Segment
X28589 N28589 N28590 Segment
X28590 N28590 N28591 Segment
X28591 N28591 N28592 Segment
X28592 N28592 N28593 Segment
X28593 N28593 N28594 Segment
X28594 N28594 N28595 Segment
X28595 N28595 N28596 Segment
X28596 N28596 N28597 Segment
X28597 N28597 N28598 Segment
X28598 N28598 N28599 Segment
X28599 N28599 N28600 Segment
X28600 N28600 N28601 Segment
X28601 N28601 N28602 Segment
X28602 N28602 N28603 Segment
X28603 N28603 N28604 Segment
X28604 N28604 N28605 Segment
X28605 N28605 N28606 Segment
X28606 N28606 N28607 Segment
X28607 N28607 N28608 Segment
X28608 N28608 N28609 Segment
X28609 N28609 N28610 Segment
X28610 N28610 N28611 Segment
X28611 N28611 N28612 Segment
X28612 N28612 N28613 Segment
X28613 N28613 N28614 Segment
X28614 N28614 N28615 Segment
X28615 N28615 N28616 Segment
X28616 N28616 N28617 Segment
X28617 N28617 N28618 Segment
X28618 N28618 N28619 Segment
X28619 N28619 N28620 Segment
X28620 N28620 N28621 Segment
X28621 N28621 N28622 Segment
X28622 N28622 N28623 Segment
X28623 N28623 N28624 Segment
X28624 N28624 N28625 Segment
X28625 N28625 N28626 Segment
X28626 N28626 N28627 Segment
X28627 N28627 N28628 Segment
X28628 N28628 N28629 Segment
X28629 N28629 N28630 Segment
X28630 N28630 N28631 Segment
X28631 N28631 N28632 Segment
X28632 N28632 N28633 Segment
X28633 N28633 N28634 Segment
X28634 N28634 N28635 Segment
X28635 N28635 N28636 Segment
X28636 N28636 N28637 Segment
X28637 N28637 N28638 Segment
X28638 N28638 N28639 Segment
X28639 N28639 N28640 Segment
X28640 N28640 N28641 Segment
X28641 N28641 N28642 Segment
X28642 N28642 N28643 Segment
X28643 N28643 N28644 Segment
X28644 N28644 N28645 Segment
X28645 N28645 N28646 Segment
X28646 N28646 N28647 Segment
X28647 N28647 N28648 Segment
X28648 N28648 N28649 Segment
X28649 N28649 N28650 Segment
X28650 N28650 N28651 Segment
X28651 N28651 N28652 Segment
X28652 N28652 N28653 Segment
X28653 N28653 N28654 Segment
X28654 N28654 N28655 Segment
X28655 N28655 N28656 Segment
X28656 N28656 N28657 Segment
X28657 N28657 N28658 Segment
X28658 N28658 N28659 Segment
X28659 N28659 N28660 Segment
X28660 N28660 N28661 Segment
X28661 N28661 N28662 Segment
X28662 N28662 N28663 Segment
X28663 N28663 N28664 Segment
X28664 N28664 N28665 Segment
X28665 N28665 N28666 Segment
X28666 N28666 N28667 Segment
X28667 N28667 N28668 Segment
X28668 N28668 N28669 Segment
X28669 N28669 N28670 Segment
X28670 N28670 N28671 Segment
X28671 N28671 N28672 Segment
X28672 N28672 N28673 Segment
X28673 N28673 N28674 Segment
X28674 N28674 N28675 Segment
X28675 N28675 N28676 Segment
X28676 N28676 N28677 Segment
X28677 N28677 N28678 Segment
X28678 N28678 N28679 Segment
X28679 N28679 N28680 Segment
X28680 N28680 N28681 Segment
X28681 N28681 N28682 Segment
X28682 N28682 N28683 Segment
X28683 N28683 N28684 Segment
X28684 N28684 N28685 Segment
X28685 N28685 N28686 Segment
X28686 N28686 N28687 Segment
X28687 N28687 N28688 Segment
X28688 N28688 N28689 Segment
X28689 N28689 N28690 Segment
X28690 N28690 N28691 Segment
X28691 N28691 N28692 Segment
X28692 N28692 N28693 Segment
X28693 N28693 N28694 Segment
X28694 N28694 N28695 Segment
X28695 N28695 N28696 Segment
X28696 N28696 N28697 Segment
X28697 N28697 N28698 Segment
X28698 N28698 N28699 Segment
X28699 N28699 N28700 Segment
X28700 N28700 N28701 Segment
X28701 N28701 N28702 Segment
X28702 N28702 N28703 Segment
X28703 N28703 N28704 Segment
X28704 N28704 N28705 Segment
X28705 N28705 N28706 Segment
X28706 N28706 N28707 Segment
X28707 N28707 N28708 Segment
X28708 N28708 N28709 Segment
X28709 N28709 N28710 Segment
X28710 N28710 N28711 Segment
X28711 N28711 N28712 Segment
X28712 N28712 N28713 Segment
X28713 N28713 N28714 Segment
X28714 N28714 N28715 Segment
X28715 N28715 N28716 Segment
X28716 N28716 N28717 Segment
X28717 N28717 N28718 Segment
X28718 N28718 N28719 Segment
X28719 N28719 N28720 Segment
X28720 N28720 N28721 Segment
X28721 N28721 N28722 Segment
X28722 N28722 N28723 Segment
X28723 N28723 N28724 Segment
X28724 N28724 N28725 Segment
X28725 N28725 N28726 Segment
X28726 N28726 N28727 Segment
X28727 N28727 N28728 Segment
X28728 N28728 N28729 Segment
X28729 N28729 N28730 Segment
X28730 N28730 N28731 Segment
X28731 N28731 N28732 Segment
X28732 N28732 N28733 Segment
X28733 N28733 N28734 Segment
X28734 N28734 N28735 Segment
X28735 N28735 N28736 Segment
X28736 N28736 N28737 Segment
X28737 N28737 N28738 Segment
X28738 N28738 N28739 Segment
X28739 N28739 N28740 Segment
X28740 N28740 N28741 Segment
X28741 N28741 N28742 Segment
X28742 N28742 N28743 Segment
X28743 N28743 N28744 Segment
X28744 N28744 N28745 Segment
X28745 N28745 N28746 Segment
X28746 N28746 N28747 Segment
X28747 N28747 N28748 Segment
X28748 N28748 N28749 Segment
X28749 N28749 N28750 Segment
X28750 N28750 N28751 Segment
X28751 N28751 N28752 Segment
X28752 N28752 N28753 Segment
X28753 N28753 N28754 Segment
X28754 N28754 N28755 Segment
X28755 N28755 N28756 Segment
X28756 N28756 N28757 Segment
X28757 N28757 N28758 Segment
X28758 N28758 N28759 Segment
X28759 N28759 N28760 Segment
X28760 N28760 N28761 Segment
X28761 N28761 N28762 Segment
X28762 N28762 N28763 Segment
X28763 N28763 N28764 Segment
X28764 N28764 N28765 Segment
X28765 N28765 N28766 Segment
X28766 N28766 N28767 Segment
X28767 N28767 N28768 Segment
X28768 N28768 N28769 Segment
X28769 N28769 N28770 Segment
X28770 N28770 N28771 Segment
X28771 N28771 N28772 Segment
X28772 N28772 N28773 Segment
X28773 N28773 N28774 Segment
X28774 N28774 N28775 Segment
X28775 N28775 N28776 Segment
X28776 N28776 N28777 Segment
X28777 N28777 N28778 Segment
X28778 N28778 N28779 Segment
X28779 N28779 N28780 Segment
X28780 N28780 N28781 Segment
X28781 N28781 N28782 Segment
X28782 N28782 N28783 Segment
X28783 N28783 N28784 Segment
X28784 N28784 N28785 Segment
X28785 N28785 N28786 Segment
X28786 N28786 N28787 Segment
X28787 N28787 N28788 Segment
X28788 N28788 N28789 Segment
X28789 N28789 N28790 Segment
X28790 N28790 N28791 Segment
X28791 N28791 N28792 Segment
X28792 N28792 N28793 Segment
X28793 N28793 N28794 Segment
X28794 N28794 N28795 Segment
X28795 N28795 N28796 Segment
X28796 N28796 N28797 Segment
X28797 N28797 N28798 Segment
X28798 N28798 N28799 Segment
X28799 N28799 N28800 Segment
X28800 N28800 N28801 Segment
X28801 N28801 N28802 Segment
X28802 N28802 N28803 Segment
X28803 N28803 N28804 Segment
X28804 N28804 N28805 Segment
X28805 N28805 N28806 Segment
X28806 N28806 N28807 Segment
X28807 N28807 N28808 Segment
X28808 N28808 N28809 Segment
X28809 N28809 N28810 Segment
X28810 N28810 N28811 Segment
X28811 N28811 N28812 Segment
X28812 N28812 N28813 Segment
X28813 N28813 N28814 Segment
X28814 N28814 N28815 Segment
X28815 N28815 N28816 Segment
X28816 N28816 N28817 Segment
X28817 N28817 N28818 Segment
X28818 N28818 N28819 Segment
X28819 N28819 N28820 Segment
X28820 N28820 N28821 Segment
X28821 N28821 N28822 Segment
X28822 N28822 N28823 Segment
X28823 N28823 N28824 Segment
X28824 N28824 N28825 Segment
X28825 N28825 N28826 Segment
X28826 N28826 N28827 Segment
X28827 N28827 N28828 Segment
X28828 N28828 N28829 Segment
X28829 N28829 N28830 Segment
X28830 N28830 N28831 Segment
X28831 N28831 N28832 Segment
X28832 N28832 N28833 Segment
X28833 N28833 N28834 Segment
X28834 N28834 N28835 Segment
X28835 N28835 N28836 Segment
X28836 N28836 N28837 Segment
X28837 N28837 N28838 Segment
X28838 N28838 N28839 Segment
X28839 N28839 N28840 Segment
X28840 N28840 N28841 Segment
X28841 N28841 N28842 Segment
X28842 N28842 N28843 Segment
X28843 N28843 N28844 Segment
X28844 N28844 N28845 Segment
X28845 N28845 N28846 Segment
X28846 N28846 N28847 Segment
X28847 N28847 N28848 Segment
X28848 N28848 N28849 Segment
X28849 N28849 N28850 Segment
X28850 N28850 N28851 Segment
X28851 N28851 N28852 Segment
X28852 N28852 N28853 Segment
X28853 N28853 N28854 Segment
X28854 N28854 N28855 Segment
X28855 N28855 N28856 Segment
X28856 N28856 N28857 Segment
X28857 N28857 N28858 Segment
X28858 N28858 N28859 Segment
X28859 N28859 N28860 Segment
X28860 N28860 N28861 Segment
X28861 N28861 N28862 Segment
X28862 N28862 N28863 Segment
X28863 N28863 N28864 Segment
X28864 N28864 N28865 Segment
X28865 N28865 N28866 Segment
X28866 N28866 N28867 Segment
X28867 N28867 N28868 Segment
X28868 N28868 N28869 Segment
X28869 N28869 N28870 Segment
X28870 N28870 N28871 Segment
X28871 N28871 N28872 Segment
X28872 N28872 N28873 Segment
X28873 N28873 N28874 Segment
X28874 N28874 N28875 Segment
X28875 N28875 N28876 Segment
X28876 N28876 N28877 Segment
X28877 N28877 N28878 Segment
X28878 N28878 N28879 Segment
X28879 N28879 N28880 Segment
X28880 N28880 N28881 Segment
X28881 N28881 N28882 Segment
X28882 N28882 N28883 Segment
X28883 N28883 N28884 Segment
X28884 N28884 N28885 Segment
X28885 N28885 N28886 Segment
X28886 N28886 N28887 Segment
X28887 N28887 N28888 Segment
X28888 N28888 N28889 Segment
X28889 N28889 N28890 Segment
X28890 N28890 N28891 Segment
X28891 N28891 N28892 Segment
X28892 N28892 N28893 Segment
X28893 N28893 N28894 Segment
X28894 N28894 N28895 Segment
X28895 N28895 N28896 Segment
X28896 N28896 N28897 Segment
X28897 N28897 N28898 Segment
X28898 N28898 N28899 Segment
X28899 N28899 N28900 Segment
X28900 N28900 N28901 Segment
X28901 N28901 N28902 Segment
X28902 N28902 N28903 Segment
X28903 N28903 N28904 Segment
X28904 N28904 N28905 Segment
X28905 N28905 N28906 Segment
X28906 N28906 N28907 Segment
X28907 N28907 N28908 Segment
X28908 N28908 N28909 Segment
X28909 N28909 N28910 Segment
X28910 N28910 N28911 Segment
X28911 N28911 N28912 Segment
X28912 N28912 N28913 Segment
X28913 N28913 N28914 Segment
X28914 N28914 N28915 Segment
X28915 N28915 N28916 Segment
X28916 N28916 N28917 Segment
X28917 N28917 N28918 Segment
X28918 N28918 N28919 Segment
X28919 N28919 N28920 Segment
X28920 N28920 N28921 Segment
X28921 N28921 N28922 Segment
X28922 N28922 N28923 Segment
X28923 N28923 N28924 Segment
X28924 N28924 N28925 Segment
X28925 N28925 N28926 Segment
X28926 N28926 N28927 Segment
X28927 N28927 N28928 Segment
X28928 N28928 N28929 Segment
X28929 N28929 N28930 Segment
X28930 N28930 N28931 Segment
X28931 N28931 N28932 Segment
X28932 N28932 N28933 Segment
X28933 N28933 N28934 Segment
X28934 N28934 N28935 Segment
X28935 N28935 N28936 Segment
X28936 N28936 N28937 Segment
X28937 N28937 N28938 Segment
X28938 N28938 N28939 Segment
X28939 N28939 N28940 Segment
X28940 N28940 N28941 Segment
X28941 N28941 N28942 Segment
X28942 N28942 N28943 Segment
X28943 N28943 N28944 Segment
X28944 N28944 N28945 Segment
X28945 N28945 N28946 Segment
X28946 N28946 N28947 Segment
X28947 N28947 N28948 Segment
X28948 N28948 N28949 Segment
X28949 N28949 N28950 Segment
X28950 N28950 N28951 Segment
X28951 N28951 N28952 Segment
X28952 N28952 N28953 Segment
X28953 N28953 N28954 Segment
X28954 N28954 N28955 Segment
X28955 N28955 N28956 Segment
X28956 N28956 N28957 Segment
X28957 N28957 N28958 Segment
X28958 N28958 N28959 Segment
X28959 N28959 N28960 Segment
X28960 N28960 N28961 Segment
X28961 N28961 N28962 Segment
X28962 N28962 N28963 Segment
X28963 N28963 N28964 Segment
X28964 N28964 N28965 Segment
X28965 N28965 N28966 Segment
X28966 N28966 N28967 Segment
X28967 N28967 N28968 Segment
X28968 N28968 N28969 Segment
X28969 N28969 N28970 Segment
X28970 N28970 N28971 Segment
X28971 N28971 N28972 Segment
X28972 N28972 N28973 Segment
X28973 N28973 N28974 Segment
X28974 N28974 N28975 Segment
X28975 N28975 N28976 Segment
X28976 N28976 N28977 Segment
X28977 N28977 N28978 Segment
X28978 N28978 N28979 Segment
X28979 N28979 N28980 Segment
X28980 N28980 N28981 Segment
X28981 N28981 N28982 Segment
X28982 N28982 N28983 Segment
X28983 N28983 N28984 Segment
X28984 N28984 N28985 Segment
X28985 N28985 N28986 Segment
X28986 N28986 N28987 Segment
X28987 N28987 N28988 Segment
X28988 N28988 N28989 Segment
X28989 N28989 N28990 Segment
X28990 N28990 N28991 Segment
X28991 N28991 N28992 Segment
X28992 N28992 N28993 Segment
X28993 N28993 N28994 Segment
X28994 N28994 N28995 Segment
X28995 N28995 N28996 Segment
X28996 N28996 N28997 Segment
X28997 N28997 N28998 Segment
X28998 N28998 N28999 Segment
X28999 N28999 N29000 Segment
X29000 N29000 N29001 Segment
X29001 N29001 N29002 Segment
X29002 N29002 N29003 Segment
X29003 N29003 N29004 Segment
X29004 N29004 N29005 Segment
X29005 N29005 N29006 Segment
X29006 N29006 N29007 Segment
X29007 N29007 N29008 Segment
X29008 N29008 N29009 Segment
X29009 N29009 N29010 Segment
X29010 N29010 N29011 Segment
X29011 N29011 N29012 Segment
X29012 N29012 N29013 Segment
X29013 N29013 N29014 Segment
X29014 N29014 N29015 Segment
X29015 N29015 N29016 Segment
X29016 N29016 N29017 Segment
X29017 N29017 N29018 Segment
X29018 N29018 N29019 Segment
X29019 N29019 N29020 Segment
X29020 N29020 N29021 Segment
X29021 N29021 N29022 Segment
X29022 N29022 N29023 Segment
X29023 N29023 N29024 Segment
X29024 N29024 N29025 Segment
X29025 N29025 N29026 Segment
X29026 N29026 N29027 Segment
X29027 N29027 N29028 Segment
X29028 N29028 N29029 Segment
X29029 N29029 N29030 Segment
X29030 N29030 N29031 Segment
X29031 N29031 N29032 Segment
X29032 N29032 N29033 Segment
X29033 N29033 N29034 Segment
X29034 N29034 N29035 Segment
X29035 N29035 N29036 Segment
X29036 N29036 N29037 Segment
X29037 N29037 N29038 Segment
X29038 N29038 N29039 Segment
X29039 N29039 N29040 Segment
X29040 N29040 N29041 Segment
X29041 N29041 N29042 Segment
X29042 N29042 N29043 Segment
X29043 N29043 N29044 Segment
X29044 N29044 N29045 Segment
X29045 N29045 N29046 Segment
X29046 N29046 N29047 Segment
X29047 N29047 N29048 Segment
X29048 N29048 N29049 Segment
X29049 N29049 N29050 Segment
X29050 N29050 N29051 Segment
X29051 N29051 N29052 Segment
X29052 N29052 N29053 Segment
X29053 N29053 N29054 Segment
X29054 N29054 N29055 Segment
X29055 N29055 N29056 Segment
X29056 N29056 N29057 Segment
X29057 N29057 N29058 Segment
X29058 N29058 N29059 Segment
X29059 N29059 N29060 Segment
X29060 N29060 N29061 Segment
X29061 N29061 N29062 Segment
X29062 N29062 N29063 Segment
X29063 N29063 N29064 Segment
X29064 N29064 N29065 Segment
X29065 N29065 N29066 Segment
X29066 N29066 N29067 Segment
X29067 N29067 N29068 Segment
X29068 N29068 N29069 Segment
X29069 N29069 N29070 Segment
X29070 N29070 N29071 Segment
X29071 N29071 N29072 Segment
X29072 N29072 N29073 Segment
X29073 N29073 N29074 Segment
X29074 N29074 N29075 Segment
X29075 N29075 N29076 Segment
X29076 N29076 N29077 Segment
X29077 N29077 N29078 Segment
X29078 N29078 N29079 Segment
X29079 N29079 N29080 Segment
X29080 N29080 N29081 Segment
X29081 N29081 N29082 Segment
X29082 N29082 N29083 Segment
X29083 N29083 N29084 Segment
X29084 N29084 N29085 Segment
X29085 N29085 N29086 Segment
X29086 N29086 N29087 Segment
X29087 N29087 N29088 Segment
X29088 N29088 N29089 Segment
X29089 N29089 N29090 Segment
X29090 N29090 N29091 Segment
X29091 N29091 N29092 Segment
X29092 N29092 N29093 Segment
X29093 N29093 N29094 Segment
X29094 N29094 N29095 Segment
X29095 N29095 N29096 Segment
X29096 N29096 N29097 Segment
X29097 N29097 N29098 Segment
X29098 N29098 N29099 Segment
X29099 N29099 N29100 Segment
X29100 N29100 N29101 Segment
X29101 N29101 N29102 Segment
X29102 N29102 N29103 Segment
X29103 N29103 N29104 Segment
X29104 N29104 N29105 Segment
X29105 N29105 N29106 Segment
X29106 N29106 N29107 Segment
X29107 N29107 N29108 Segment
X29108 N29108 N29109 Segment
X29109 N29109 N29110 Segment
X29110 N29110 N29111 Segment
X29111 N29111 N29112 Segment
X29112 N29112 N29113 Segment
X29113 N29113 N29114 Segment
X29114 N29114 N29115 Segment
X29115 N29115 N29116 Segment
X29116 N29116 N29117 Segment
X29117 N29117 N29118 Segment
X29118 N29118 N29119 Segment
X29119 N29119 N29120 Segment
X29120 N29120 N29121 Segment
X29121 N29121 N29122 Segment
X29122 N29122 N29123 Segment
X29123 N29123 N29124 Segment
X29124 N29124 N29125 Segment
X29125 N29125 N29126 Segment
X29126 N29126 N29127 Segment
X29127 N29127 N29128 Segment
X29128 N29128 N29129 Segment
X29129 N29129 N29130 Segment
X29130 N29130 N29131 Segment
X29131 N29131 N29132 Segment
X29132 N29132 N29133 Segment
X29133 N29133 N29134 Segment
X29134 N29134 N29135 Segment
X29135 N29135 N29136 Segment
X29136 N29136 N29137 Segment
X29137 N29137 N29138 Segment
X29138 N29138 N29139 Segment
X29139 N29139 N29140 Segment
X29140 N29140 N29141 Segment
X29141 N29141 N29142 Segment
X29142 N29142 N29143 Segment
X29143 N29143 N29144 Segment
X29144 N29144 N29145 Segment
X29145 N29145 N29146 Segment
X29146 N29146 N29147 Segment
X29147 N29147 N29148 Segment
X29148 N29148 N29149 Segment
X29149 N29149 N29150 Segment
X29150 N29150 N29151 Segment
X29151 N29151 N29152 Segment
X29152 N29152 N29153 Segment
X29153 N29153 N29154 Segment
X29154 N29154 N29155 Segment
X29155 N29155 N29156 Segment
X29156 N29156 N29157 Segment
X29157 N29157 N29158 Segment
X29158 N29158 N29159 Segment
X29159 N29159 N29160 Segment
X29160 N29160 N29161 Segment
X29161 N29161 N29162 Segment
X29162 N29162 N29163 Segment
X29163 N29163 N29164 Segment
X29164 N29164 N29165 Segment
X29165 N29165 N29166 Segment
X29166 N29166 N29167 Segment
X29167 N29167 N29168 Segment
X29168 N29168 N29169 Segment
X29169 N29169 N29170 Segment
X29170 N29170 N29171 Segment
X29171 N29171 N29172 Segment
X29172 N29172 N29173 Segment
X29173 N29173 N29174 Segment
X29174 N29174 N29175 Segment
X29175 N29175 N29176 Segment
X29176 N29176 N29177 Segment
X29177 N29177 N29178 Segment
X29178 N29178 N29179 Segment
X29179 N29179 N29180 Segment
X29180 N29180 N29181 Segment
X29181 N29181 N29182 Segment
X29182 N29182 N29183 Segment
X29183 N29183 N29184 Segment
X29184 N29184 N29185 Segment
X29185 N29185 N29186 Segment
X29186 N29186 N29187 Segment
X29187 N29187 N29188 Segment
X29188 N29188 N29189 Segment
X29189 N29189 N29190 Segment
X29190 N29190 N29191 Segment
X29191 N29191 N29192 Segment
X29192 N29192 N29193 Segment
X29193 N29193 N29194 Segment
X29194 N29194 N29195 Segment
X29195 N29195 N29196 Segment
X29196 N29196 N29197 Segment
X29197 N29197 N29198 Segment
X29198 N29198 N29199 Segment
X29199 N29199 N29200 Segment
X29200 N29200 N29201 Segment
X29201 N29201 N29202 Segment
X29202 N29202 N29203 Segment
X29203 N29203 N29204 Segment
X29204 N29204 N29205 Segment
X29205 N29205 N29206 Segment
X29206 N29206 N29207 Segment
X29207 N29207 N29208 Segment
X29208 N29208 N29209 Segment
X29209 N29209 N29210 Segment
X29210 N29210 N29211 Segment
X29211 N29211 N29212 Segment
X29212 N29212 N29213 Segment
X29213 N29213 N29214 Segment
X29214 N29214 N29215 Segment
X29215 N29215 N29216 Segment
X29216 N29216 N29217 Segment
X29217 N29217 N29218 Segment
X29218 N29218 N29219 Segment
X29219 N29219 N29220 Segment
X29220 N29220 N29221 Segment
X29221 N29221 N29222 Segment
X29222 N29222 N29223 Segment
X29223 N29223 N29224 Segment
X29224 N29224 N29225 Segment
X29225 N29225 N29226 Segment
X29226 N29226 N29227 Segment
X29227 N29227 N29228 Segment
X29228 N29228 N29229 Segment
X29229 N29229 N29230 Segment
X29230 N29230 N29231 Segment
X29231 N29231 N29232 Segment
X29232 N29232 N29233 Segment
X29233 N29233 N29234 Segment
X29234 N29234 N29235 Segment
X29235 N29235 N29236 Segment
X29236 N29236 N29237 Segment
X29237 N29237 N29238 Segment
X29238 N29238 N29239 Segment
X29239 N29239 N29240 Segment
X29240 N29240 N29241 Segment
X29241 N29241 N29242 Segment
X29242 N29242 N29243 Segment
X29243 N29243 N29244 Segment
X29244 N29244 N29245 Segment
X29245 N29245 N29246 Segment
X29246 N29246 N29247 Segment
X29247 N29247 N29248 Segment
X29248 N29248 N29249 Segment
X29249 N29249 N29250 Segment
X29250 N29250 N29251 Segment
X29251 N29251 N29252 Segment
X29252 N29252 N29253 Segment
X29253 N29253 N29254 Segment
X29254 N29254 N29255 Segment
X29255 N29255 N29256 Segment
X29256 N29256 N29257 Segment
X29257 N29257 N29258 Segment
X29258 N29258 N29259 Segment
X29259 N29259 N29260 Segment
X29260 N29260 N29261 Segment
X29261 N29261 N29262 Segment
X29262 N29262 N29263 Segment
X29263 N29263 N29264 Segment
X29264 N29264 N29265 Segment
X29265 N29265 N29266 Segment
X29266 N29266 N29267 Segment
X29267 N29267 N29268 Segment
X29268 N29268 N29269 Segment
X29269 N29269 N29270 Segment
X29270 N29270 N29271 Segment
X29271 N29271 N29272 Segment
X29272 N29272 N29273 Segment
X29273 N29273 N29274 Segment
X29274 N29274 N29275 Segment
X29275 N29275 N29276 Segment
X29276 N29276 N29277 Segment
X29277 N29277 N29278 Segment
X29278 N29278 N29279 Segment
X29279 N29279 N29280 Segment
X29280 N29280 N29281 Segment
X29281 N29281 N29282 Segment
X29282 N29282 N29283 Segment
X29283 N29283 N29284 Segment
X29284 N29284 N29285 Segment
X29285 N29285 N29286 Segment
X29286 N29286 N29287 Segment
X29287 N29287 N29288 Segment
X29288 N29288 N29289 Segment
X29289 N29289 N29290 Segment
X29290 N29290 N29291 Segment
X29291 N29291 N29292 Segment
X29292 N29292 N29293 Segment
X29293 N29293 N29294 Segment
X29294 N29294 N29295 Segment
X29295 N29295 N29296 Segment
X29296 N29296 N29297 Segment
X29297 N29297 N29298 Segment
X29298 N29298 N29299 Segment
X29299 N29299 N29300 Segment
X29300 N29300 N29301 Segment
X29301 N29301 N29302 Segment
X29302 N29302 N29303 Segment
X29303 N29303 N29304 Segment
X29304 N29304 N29305 Segment
X29305 N29305 N29306 Segment
X29306 N29306 N29307 Segment
X29307 N29307 N29308 Segment
X29308 N29308 N29309 Segment
X29309 N29309 N29310 Segment
X29310 N29310 N29311 Segment
X29311 N29311 N29312 Segment
X29312 N29312 N29313 Segment
X29313 N29313 N29314 Segment
X29314 N29314 N29315 Segment
X29315 N29315 N29316 Segment
X29316 N29316 N29317 Segment
X29317 N29317 N29318 Segment
X29318 N29318 N29319 Segment
X29319 N29319 N29320 Segment
X29320 N29320 N29321 Segment
X29321 N29321 N29322 Segment
X29322 N29322 N29323 Segment
X29323 N29323 N29324 Segment
X29324 N29324 N29325 Segment
X29325 N29325 N29326 Segment
X29326 N29326 N29327 Segment
X29327 N29327 N29328 Segment
X29328 N29328 N29329 Segment
X29329 N29329 N29330 Segment
X29330 N29330 N29331 Segment
X29331 N29331 N29332 Segment
X29332 N29332 N29333 Segment
X29333 N29333 N29334 Segment
X29334 N29334 N29335 Segment
X29335 N29335 N29336 Segment
X29336 N29336 N29337 Segment
X29337 N29337 N29338 Segment
X29338 N29338 N29339 Segment
X29339 N29339 N29340 Segment
X29340 N29340 N29341 Segment
X29341 N29341 N29342 Segment
X29342 N29342 N29343 Segment
X29343 N29343 N29344 Segment
X29344 N29344 N29345 Segment
X29345 N29345 N29346 Segment
X29346 N29346 N29347 Segment
X29347 N29347 N29348 Segment
X29348 N29348 N29349 Segment
X29349 N29349 N29350 Segment
X29350 N29350 N29351 Segment
X29351 N29351 N29352 Segment
X29352 N29352 N29353 Segment
X29353 N29353 N29354 Segment
X29354 N29354 N29355 Segment
X29355 N29355 N29356 Segment
X29356 N29356 N29357 Segment
X29357 N29357 N29358 Segment
X29358 N29358 N29359 Segment
X29359 N29359 N29360 Segment
X29360 N29360 N29361 Segment
X29361 N29361 N29362 Segment
X29362 N29362 N29363 Segment
X29363 N29363 N29364 Segment
X29364 N29364 N29365 Segment
X29365 N29365 N29366 Segment
X29366 N29366 N29367 Segment
X29367 N29367 N29368 Segment
X29368 N29368 N29369 Segment
X29369 N29369 N29370 Segment
X29370 N29370 N29371 Segment
X29371 N29371 N29372 Segment
X29372 N29372 N29373 Segment
X29373 N29373 N29374 Segment
X29374 N29374 N29375 Segment
X29375 N29375 N29376 Segment
X29376 N29376 N29377 Segment
X29377 N29377 N29378 Segment
X29378 N29378 N29379 Segment
X29379 N29379 N29380 Segment
X29380 N29380 N29381 Segment
X29381 N29381 N29382 Segment
X29382 N29382 N29383 Segment
X29383 N29383 N29384 Segment
X29384 N29384 N29385 Segment
X29385 N29385 N29386 Segment
X29386 N29386 N29387 Segment
X29387 N29387 N29388 Segment
X29388 N29388 N29389 Segment
X29389 N29389 N29390 Segment
X29390 N29390 N29391 Segment
X29391 N29391 N29392 Segment
X29392 N29392 N29393 Segment
X29393 N29393 N29394 Segment
X29394 N29394 N29395 Segment
X29395 N29395 N29396 Segment
X29396 N29396 N29397 Segment
X29397 N29397 N29398 Segment
X29398 N29398 N29399 Segment
X29399 N29399 N29400 Segment
X29400 N29400 N29401 Segment
X29401 N29401 N29402 Segment
X29402 N29402 N29403 Segment
X29403 N29403 N29404 Segment
X29404 N29404 N29405 Segment
X29405 N29405 N29406 Segment
X29406 N29406 N29407 Segment
X29407 N29407 N29408 Segment
X29408 N29408 N29409 Segment
X29409 N29409 N29410 Segment
X29410 N29410 N29411 Segment
X29411 N29411 N29412 Segment
X29412 N29412 N29413 Segment
X29413 N29413 N29414 Segment
X29414 N29414 N29415 Segment
X29415 N29415 N29416 Segment
X29416 N29416 N29417 Segment
X29417 N29417 N29418 Segment
X29418 N29418 N29419 Segment
X29419 N29419 N29420 Segment
X29420 N29420 N29421 Segment
X29421 N29421 N29422 Segment
X29422 N29422 N29423 Segment
X29423 N29423 N29424 Segment
X29424 N29424 N29425 Segment
X29425 N29425 N29426 Segment
X29426 N29426 N29427 Segment
X29427 N29427 N29428 Segment
X29428 N29428 N29429 Segment
X29429 N29429 N29430 Segment
X29430 N29430 N29431 Segment
X29431 N29431 N29432 Segment
X29432 N29432 N29433 Segment
X29433 N29433 N29434 Segment
X29434 N29434 N29435 Segment
X29435 N29435 N29436 Segment
X29436 N29436 N29437 Segment
X29437 N29437 N29438 Segment
X29438 N29438 N29439 Segment
X29439 N29439 N29440 Segment
X29440 N29440 N29441 Segment
X29441 N29441 N29442 Segment
X29442 N29442 N29443 Segment
X29443 N29443 N29444 Segment
X29444 N29444 N29445 Segment
X29445 N29445 N29446 Segment
X29446 N29446 N29447 Segment
X29447 N29447 N29448 Segment
X29448 N29448 N29449 Segment
X29449 N29449 N29450 Segment
X29450 N29450 N29451 Segment
X29451 N29451 N29452 Segment
X29452 N29452 N29453 Segment
X29453 N29453 N29454 Segment
X29454 N29454 N29455 Segment
X29455 N29455 N29456 Segment
X29456 N29456 N29457 Segment
X29457 N29457 N29458 Segment
X29458 N29458 N29459 Segment
X29459 N29459 N29460 Segment
X29460 N29460 N29461 Segment
X29461 N29461 N29462 Segment
X29462 N29462 N29463 Segment
X29463 N29463 N29464 Segment
X29464 N29464 N29465 Segment
X29465 N29465 N29466 Segment
X29466 N29466 N29467 Segment
X29467 N29467 N29468 Segment
X29468 N29468 N29469 Segment
X29469 N29469 N29470 Segment
X29470 N29470 N29471 Segment
X29471 N29471 N29472 Segment
X29472 N29472 N29473 Segment
X29473 N29473 N29474 Segment
X29474 N29474 N29475 Segment
X29475 N29475 N29476 Segment
X29476 N29476 N29477 Segment
X29477 N29477 N29478 Segment
X29478 N29478 N29479 Segment
X29479 N29479 N29480 Segment
X29480 N29480 N29481 Segment
X29481 N29481 N29482 Segment
X29482 N29482 N29483 Segment
X29483 N29483 N29484 Segment
X29484 N29484 N29485 Segment
X29485 N29485 N29486 Segment
X29486 N29486 N29487 Segment
X29487 N29487 N29488 Segment
X29488 N29488 N29489 Segment
X29489 N29489 N29490 Segment
X29490 N29490 N29491 Segment
X29491 N29491 N29492 Segment
X29492 N29492 N29493 Segment
X29493 N29493 N29494 Segment
X29494 N29494 N29495 Segment
X29495 N29495 N29496 Segment
X29496 N29496 N29497 Segment
X29497 N29497 N29498 Segment
X29498 N29498 N29499 Segment
X29499 N29499 N29500 Segment
X29500 N29500 N29501 Segment
X29501 N29501 N29502 Segment
X29502 N29502 N29503 Segment
X29503 N29503 N29504 Segment
X29504 N29504 N29505 Segment
X29505 N29505 N29506 Segment
X29506 N29506 N29507 Segment
X29507 N29507 N29508 Segment
X29508 N29508 N29509 Segment
X29509 N29509 N29510 Segment
X29510 N29510 N29511 Segment
X29511 N29511 N29512 Segment
X29512 N29512 N29513 Segment
X29513 N29513 N29514 Segment
X29514 N29514 N29515 Segment
X29515 N29515 N29516 Segment
X29516 N29516 N29517 Segment
X29517 N29517 N29518 Segment
X29518 N29518 N29519 Segment
X29519 N29519 N29520 Segment
X29520 N29520 N29521 Segment
X29521 N29521 N29522 Segment
X29522 N29522 N29523 Segment
X29523 N29523 N29524 Segment
X29524 N29524 N29525 Segment
X29525 N29525 N29526 Segment
X29526 N29526 N29527 Segment
X29527 N29527 N29528 Segment
X29528 N29528 N29529 Segment
X29529 N29529 N29530 Segment
X29530 N29530 N29531 Segment
X29531 N29531 N29532 Segment
X29532 N29532 N29533 Segment
X29533 N29533 N29534 Segment
X29534 N29534 N29535 Segment
X29535 N29535 N29536 Segment
X29536 N29536 N29537 Segment
X29537 N29537 N29538 Segment
X29538 N29538 N29539 Segment
X29539 N29539 N29540 Segment
X29540 N29540 N29541 Segment
X29541 N29541 N29542 Segment
X29542 N29542 N29543 Segment
X29543 N29543 N29544 Segment
X29544 N29544 N29545 Segment
X29545 N29545 N29546 Segment
X29546 N29546 N29547 Segment
X29547 N29547 N29548 Segment
X29548 N29548 N29549 Segment
X29549 N29549 N29550 Segment
X29550 N29550 N29551 Segment
X29551 N29551 N29552 Segment
X29552 N29552 N29553 Segment
X29553 N29553 N29554 Segment
X29554 N29554 N29555 Segment
X29555 N29555 N29556 Segment
X29556 N29556 N29557 Segment
X29557 N29557 N29558 Segment
X29558 N29558 N29559 Segment
X29559 N29559 N29560 Segment
X29560 N29560 N29561 Segment
X29561 N29561 N29562 Segment
X29562 N29562 N29563 Segment
X29563 N29563 N29564 Segment
X29564 N29564 N29565 Segment
X29565 N29565 N29566 Segment
X29566 N29566 N29567 Segment
X29567 N29567 N29568 Segment
X29568 N29568 N29569 Segment
X29569 N29569 N29570 Segment
X29570 N29570 N29571 Segment
X29571 N29571 N29572 Segment
X29572 N29572 N29573 Segment
X29573 N29573 N29574 Segment
X29574 N29574 N29575 Segment
X29575 N29575 N29576 Segment
X29576 N29576 N29577 Segment
X29577 N29577 N29578 Segment
X29578 N29578 N29579 Segment
X29579 N29579 N29580 Segment
X29580 N29580 N29581 Segment
X29581 N29581 N29582 Segment
X29582 N29582 N29583 Segment
X29583 N29583 N29584 Segment
X29584 N29584 N29585 Segment
X29585 N29585 N29586 Segment
X29586 N29586 N29587 Segment
X29587 N29587 N29588 Segment
X29588 N29588 N29589 Segment
X29589 N29589 N29590 Segment
X29590 N29590 N29591 Segment
X29591 N29591 N29592 Segment
X29592 N29592 N29593 Segment
X29593 N29593 N29594 Segment
X29594 N29594 N29595 Segment
X29595 N29595 N29596 Segment
X29596 N29596 N29597 Segment
X29597 N29597 N29598 Segment
X29598 N29598 N29599 Segment
X29599 N29599 N29600 Segment
X29600 N29600 N29601 Segment
X29601 N29601 N29602 Segment
X29602 N29602 N29603 Segment
X29603 N29603 N29604 Segment
X29604 N29604 N29605 Segment
X29605 N29605 N29606 Segment
X29606 N29606 N29607 Segment
X29607 N29607 N29608 Segment
X29608 N29608 N29609 Segment
X29609 N29609 N29610 Segment
X29610 N29610 N29611 Segment
X29611 N29611 N29612 Segment
X29612 N29612 N29613 Segment
X29613 N29613 N29614 Segment
X29614 N29614 N29615 Segment
X29615 N29615 N29616 Segment
X29616 N29616 N29617 Segment
X29617 N29617 N29618 Segment
X29618 N29618 N29619 Segment
X29619 N29619 N29620 Segment
X29620 N29620 N29621 Segment
X29621 N29621 N29622 Segment
X29622 N29622 N29623 Segment
X29623 N29623 N29624 Segment
X29624 N29624 N29625 Segment
X29625 N29625 N29626 Segment
X29626 N29626 N29627 Segment
X29627 N29627 N29628 Segment
X29628 N29628 N29629 Segment
X29629 N29629 N29630 Segment
X29630 N29630 N29631 Segment
X29631 N29631 N29632 Segment
X29632 N29632 N29633 Segment
X29633 N29633 N29634 Segment
X29634 N29634 N29635 Segment
X29635 N29635 N29636 Segment
X29636 N29636 N29637 Segment
X29637 N29637 N29638 Segment
X29638 N29638 N29639 Segment
X29639 N29639 N29640 Segment
X29640 N29640 N29641 Segment
X29641 N29641 N29642 Segment
X29642 N29642 N29643 Segment
X29643 N29643 N29644 Segment
X29644 N29644 N29645 Segment
X29645 N29645 N29646 Segment
X29646 N29646 N29647 Segment
X29647 N29647 N29648 Segment
X29648 N29648 N29649 Segment
X29649 N29649 N29650 Segment
X29650 N29650 N29651 Segment
X29651 N29651 N29652 Segment
X29652 N29652 N29653 Segment
X29653 N29653 N29654 Segment
X29654 N29654 N29655 Segment
X29655 N29655 N29656 Segment
X29656 N29656 N29657 Segment
X29657 N29657 N29658 Segment
X29658 N29658 N29659 Segment
X29659 N29659 N29660 Segment
X29660 N29660 N29661 Segment
X29661 N29661 N29662 Segment
X29662 N29662 N29663 Segment
X29663 N29663 N29664 Segment
X29664 N29664 N29665 Segment
X29665 N29665 N29666 Segment
X29666 N29666 N29667 Segment
X29667 N29667 N29668 Segment
X29668 N29668 N29669 Segment
X29669 N29669 N29670 Segment
X29670 N29670 N29671 Segment
X29671 N29671 N29672 Segment
X29672 N29672 N29673 Segment
X29673 N29673 N29674 Segment
X29674 N29674 N29675 Segment
X29675 N29675 N29676 Segment
X29676 N29676 N29677 Segment
X29677 N29677 N29678 Segment
X29678 N29678 N29679 Segment
X29679 N29679 N29680 Segment
X29680 N29680 N29681 Segment
X29681 N29681 N29682 Segment
X29682 N29682 N29683 Segment
X29683 N29683 N29684 Segment
X29684 N29684 N29685 Segment
X29685 N29685 N29686 Segment
X29686 N29686 N29687 Segment
X29687 N29687 N29688 Segment
X29688 N29688 N29689 Segment
X29689 N29689 N29690 Segment
X29690 N29690 N29691 Segment
X29691 N29691 N29692 Segment
X29692 N29692 N29693 Segment
X29693 N29693 N29694 Segment
X29694 N29694 N29695 Segment
X29695 N29695 N29696 Segment
X29696 N29696 N29697 Segment
X29697 N29697 N29698 Segment
X29698 N29698 N29699 Segment
X29699 N29699 N29700 Segment
X29700 N29700 N29701 Segment
X29701 N29701 N29702 Segment
X29702 N29702 N29703 Segment
X29703 N29703 N29704 Segment
X29704 N29704 N29705 Segment
X29705 N29705 N29706 Segment
X29706 N29706 N29707 Segment
X29707 N29707 N29708 Segment
X29708 N29708 N29709 Segment
X29709 N29709 N29710 Segment
X29710 N29710 N29711 Segment
X29711 N29711 N29712 Segment
X29712 N29712 N29713 Segment
X29713 N29713 N29714 Segment
X29714 N29714 N29715 Segment
X29715 N29715 N29716 Segment
X29716 N29716 N29717 Segment
X29717 N29717 N29718 Segment
X29718 N29718 N29719 Segment
X29719 N29719 N29720 Segment
X29720 N29720 N29721 Segment
X29721 N29721 N29722 Segment
X29722 N29722 N29723 Segment
X29723 N29723 N29724 Segment
X29724 N29724 N29725 Segment
X29725 N29725 N29726 Segment
X29726 N29726 N29727 Segment
X29727 N29727 N29728 Segment
X29728 N29728 N29729 Segment
X29729 N29729 N29730 Segment
X29730 N29730 N29731 Segment
X29731 N29731 N29732 Segment
X29732 N29732 N29733 Segment
X29733 N29733 N29734 Segment
X29734 N29734 N29735 Segment
X29735 N29735 N29736 Segment
X29736 N29736 N29737 Segment
X29737 N29737 N29738 Segment
X29738 N29738 N29739 Segment
X29739 N29739 N29740 Segment
X29740 N29740 N29741 Segment
X29741 N29741 N29742 Segment
X29742 N29742 N29743 Segment
X29743 N29743 N29744 Segment
X29744 N29744 N29745 Segment
X29745 N29745 N29746 Segment
X29746 N29746 N29747 Segment
X29747 N29747 N29748 Segment
X29748 N29748 N29749 Segment
X29749 N29749 N29750 Segment
X29750 N29750 N29751 Segment
X29751 N29751 N29752 Segment
X29752 N29752 N29753 Segment
X29753 N29753 N29754 Segment
X29754 N29754 N29755 Segment
X29755 N29755 N29756 Segment
X29756 N29756 N29757 Segment
X29757 N29757 N29758 Segment
X29758 N29758 N29759 Segment
X29759 N29759 N29760 Segment
X29760 N29760 N29761 Segment
X29761 N29761 N29762 Segment
X29762 N29762 N29763 Segment
X29763 N29763 N29764 Segment
X29764 N29764 N29765 Segment
X29765 N29765 N29766 Segment
X29766 N29766 N29767 Segment
X29767 N29767 N29768 Segment
X29768 N29768 N29769 Segment
X29769 N29769 N29770 Segment
X29770 N29770 N29771 Segment
X29771 N29771 N29772 Segment
X29772 N29772 N29773 Segment
X29773 N29773 N29774 Segment
X29774 N29774 N29775 Segment
X29775 N29775 N29776 Segment
X29776 N29776 N29777 Segment
X29777 N29777 N29778 Segment
X29778 N29778 N29779 Segment
X29779 N29779 N29780 Segment
X29780 N29780 N29781 Segment
X29781 N29781 N29782 Segment
X29782 N29782 N29783 Segment
X29783 N29783 N29784 Segment
X29784 N29784 N29785 Segment
X29785 N29785 N29786 Segment
X29786 N29786 N29787 Segment
X29787 N29787 N29788 Segment
X29788 N29788 N29789 Segment
X29789 N29789 N29790 Segment
X29790 N29790 N29791 Segment
X29791 N29791 N29792 Segment
X29792 N29792 N29793 Segment
X29793 N29793 N29794 Segment
X29794 N29794 N29795 Segment
X29795 N29795 N29796 Segment
X29796 N29796 N29797 Segment
X29797 N29797 N29798 Segment
X29798 N29798 N29799 Segment
X29799 N29799 N29800 Segment
X29800 N29800 N29801 Segment
X29801 N29801 N29802 Segment
X29802 N29802 N29803 Segment
X29803 N29803 N29804 Segment
X29804 N29804 N29805 Segment
X29805 N29805 N29806 Segment
X29806 N29806 N29807 Segment
X29807 N29807 N29808 Segment
X29808 N29808 N29809 Segment
X29809 N29809 N29810 Segment
X29810 N29810 N29811 Segment
X29811 N29811 N29812 Segment
X29812 N29812 N29813 Segment
X29813 N29813 N29814 Segment
X29814 N29814 N29815 Segment
X29815 N29815 N29816 Segment
X29816 N29816 N29817 Segment
X29817 N29817 N29818 Segment
X29818 N29818 N29819 Segment
X29819 N29819 N29820 Segment
X29820 N29820 N29821 Segment
X29821 N29821 N29822 Segment
X29822 N29822 N29823 Segment
X29823 N29823 N29824 Segment
X29824 N29824 N29825 Segment
X29825 N29825 N29826 Segment
X29826 N29826 N29827 Segment
X29827 N29827 N29828 Segment
X29828 N29828 N29829 Segment
X29829 N29829 N29830 Segment
X29830 N29830 N29831 Segment
X29831 N29831 N29832 Segment
X29832 N29832 N29833 Segment
X29833 N29833 N29834 Segment
X29834 N29834 N29835 Segment
X29835 N29835 N29836 Segment
X29836 N29836 N29837 Segment
X29837 N29837 N29838 Segment
X29838 N29838 N29839 Segment
X29839 N29839 N29840 Segment
X29840 N29840 N29841 Segment
X29841 N29841 N29842 Segment
X29842 N29842 N29843 Segment
X29843 N29843 N29844 Segment
X29844 N29844 N29845 Segment
X29845 N29845 N29846 Segment
X29846 N29846 N29847 Segment
X29847 N29847 N29848 Segment
X29848 N29848 N29849 Segment
X29849 N29849 N29850 Segment
X29850 N29850 N29851 Segment
X29851 N29851 N29852 Segment
X29852 N29852 N29853 Segment
X29853 N29853 N29854 Segment
X29854 N29854 N29855 Segment
X29855 N29855 N29856 Segment
X29856 N29856 N29857 Segment
X29857 N29857 N29858 Segment
X29858 N29858 N29859 Segment
X29859 N29859 N29860 Segment
X29860 N29860 N29861 Segment
X29861 N29861 N29862 Segment
X29862 N29862 N29863 Segment
X29863 N29863 N29864 Segment
X29864 N29864 N29865 Segment
X29865 N29865 N29866 Segment
X29866 N29866 N29867 Segment
X29867 N29867 N29868 Segment
X29868 N29868 N29869 Segment
X29869 N29869 N29870 Segment
X29870 N29870 N29871 Segment
X29871 N29871 N29872 Segment
X29872 N29872 N29873 Segment
X29873 N29873 N29874 Segment
X29874 N29874 N29875 Segment
X29875 N29875 N29876 Segment
X29876 N29876 N29877 Segment
X29877 N29877 N29878 Segment
X29878 N29878 N29879 Segment
X29879 N29879 N29880 Segment
X29880 N29880 N29881 Segment
X29881 N29881 N29882 Segment
X29882 N29882 N29883 Segment
X29883 N29883 N29884 Segment
X29884 N29884 N29885 Segment
X29885 N29885 N29886 Segment
X29886 N29886 N29887 Segment
X29887 N29887 N29888 Segment
X29888 N29888 N29889 Segment
X29889 N29889 N29890 Segment
X29890 N29890 N29891 Segment
X29891 N29891 N29892 Segment
X29892 N29892 N29893 Segment
X29893 N29893 N29894 Segment
X29894 N29894 N29895 Segment
X29895 N29895 N29896 Segment
X29896 N29896 N29897 Segment
X29897 N29897 N29898 Segment
X29898 N29898 N29899 Segment
X29899 N29899 N29900 Segment
X29900 N29900 N29901 Segment
X29901 N29901 N29902 Segment
X29902 N29902 N29903 Segment
X29903 N29903 N29904 Segment
X29904 N29904 N29905 Segment
X29905 N29905 N29906 Segment
X29906 N29906 N29907 Segment
X29907 N29907 N29908 Segment
X29908 N29908 N29909 Segment
X29909 N29909 N29910 Segment
X29910 N29910 N29911 Segment
X29911 N29911 N29912 Segment
X29912 N29912 N29913 Segment
X29913 N29913 N29914 Segment
X29914 N29914 N29915 Segment
X29915 N29915 N29916 Segment
X29916 N29916 N29917 Segment
X29917 N29917 N29918 Segment
X29918 N29918 N29919 Segment
X29919 N29919 N29920 Segment
X29920 N29920 N29921 Segment
X29921 N29921 N29922 Segment
X29922 N29922 N29923 Segment
X29923 N29923 N29924 Segment
X29924 N29924 N29925 Segment
X29925 N29925 N29926 Segment
X29926 N29926 N29927 Segment
X29927 N29927 N29928 Segment
X29928 N29928 N29929 Segment
X29929 N29929 N29930 Segment
X29930 N29930 N29931 Segment
X29931 N29931 N29932 Segment
X29932 N29932 N29933 Segment
X29933 N29933 N29934 Segment
X29934 N29934 N29935 Segment
X29935 N29935 N29936 Segment
X29936 N29936 N29937 Segment
X29937 N29937 N29938 Segment
X29938 N29938 N29939 Segment
X29939 N29939 N29940 Segment
X29940 N29940 N29941 Segment
X29941 N29941 N29942 Segment
X29942 N29942 N29943 Segment
X29943 N29943 N29944 Segment
X29944 N29944 N29945 Segment
X29945 N29945 N29946 Segment
X29946 N29946 N29947 Segment
X29947 N29947 N29948 Segment
X29948 N29948 N29949 Segment
X29949 N29949 N29950 Segment
X29950 N29950 N29951 Segment
X29951 N29951 N29952 Segment
X29952 N29952 N29953 Segment
X29953 N29953 N29954 Segment
X29954 N29954 N29955 Segment
X29955 N29955 N29956 Segment
X29956 N29956 N29957 Segment
X29957 N29957 N29958 Segment
X29958 N29958 N29959 Segment
X29959 N29959 N29960 Segment
X29960 N29960 N29961 Segment
X29961 N29961 N29962 Segment
X29962 N29962 N29963 Segment
X29963 N29963 N29964 Segment
X29964 N29964 N29965 Segment
X29965 N29965 N29966 Segment
X29966 N29966 N29967 Segment
X29967 N29967 N29968 Segment
X29968 N29968 N29969 Segment
X29969 N29969 N29970 Segment
X29970 N29970 N29971 Segment
X29971 N29971 N29972 Segment
X29972 N29972 N29973 Segment
X29973 N29973 N29974 Segment
X29974 N29974 N29975 Segment
X29975 N29975 N29976 Segment
X29976 N29976 N29977 Segment
X29977 N29977 N29978 Segment
X29978 N29978 N29979 Segment
X29979 N29979 N29980 Segment
X29980 N29980 N29981 Segment
X29981 N29981 N29982 Segment
X29982 N29982 N29983 Segment
X29983 N29983 N29984 Segment
X29984 N29984 N29985 Segment
X29985 N29985 N29986 Segment
X29986 N29986 N29987 Segment
X29987 N29987 N29988 Segment
X29988 N29988 N29989 Segment
X29989 N29989 N29990 Segment
X29990 N29990 N29991 Segment
X29991 N29991 N29992 Segment
X29992 N29992 N29993 Segment
X29993 N29993 N29994 Segment
X29994 N29994 N29995 Segment
X29995 N29995 N29996 Segment
X29996 N29996 N29997 Segment
X29997 N29997 N29998 Segment
X29998 N29998 N29999 Segment
X29999 N29999 N30000 Segment
X30000 N30000 N30001 Segment
X30001 N30001 N30002 Segment
X30002 N30002 N30003 Segment
X30003 N30003 N30004 Segment
X30004 N30004 N30005 Segment
X30005 N30005 N30006 Segment
X30006 N30006 N30007 Segment
X30007 N30007 N30008 Segment
X30008 N30008 N30009 Segment
X30009 N30009 N30010 Segment
X30010 N30010 N30011 Segment
X30011 N30011 N30012 Segment
X30012 N30012 N30013 Segment
X30013 N30013 N30014 Segment
X30014 N30014 N30015 Segment
X30015 N30015 N30016 Segment
X30016 N30016 N30017 Segment
X30017 N30017 N30018 Segment
X30018 N30018 N30019 Segment
X30019 N30019 N30020 Segment
X30020 N30020 N30021 Segment
X30021 N30021 N30022 Segment
X30022 N30022 N30023 Segment
X30023 N30023 N30024 Segment
X30024 N30024 N30025 Segment
X30025 N30025 N30026 Segment
X30026 N30026 N30027 Segment
X30027 N30027 N30028 Segment
X30028 N30028 N30029 Segment
X30029 N30029 N30030 Segment
X30030 N30030 N30031 Segment
X30031 N30031 N30032 Segment
X30032 N30032 N30033 Segment
X30033 N30033 N30034 Segment
X30034 N30034 N30035 Segment
X30035 N30035 N30036 Segment
X30036 N30036 N30037 Segment
X30037 N30037 N30038 Segment
X30038 N30038 N30039 Segment
X30039 N30039 N30040 Segment
X30040 N30040 N30041 Segment
X30041 N30041 N30042 Segment
X30042 N30042 N30043 Segment
X30043 N30043 N30044 Segment
X30044 N30044 N30045 Segment
X30045 N30045 N30046 Segment
X30046 N30046 N30047 Segment
X30047 N30047 N30048 Segment
X30048 N30048 N30049 Segment
X30049 N30049 N30050 Segment
X30050 N30050 N30051 Segment
X30051 N30051 N30052 Segment
X30052 N30052 N30053 Segment
X30053 N30053 N30054 Segment
X30054 N30054 N30055 Segment
X30055 N30055 N30056 Segment
X30056 N30056 N30057 Segment
X30057 N30057 N30058 Segment
X30058 N30058 N30059 Segment
X30059 N30059 N30060 Segment
X30060 N30060 N30061 Segment
X30061 N30061 N30062 Segment
X30062 N30062 N30063 Segment
X30063 N30063 N30064 Segment
X30064 N30064 N30065 Segment
X30065 N30065 N30066 Segment
X30066 N30066 N30067 Segment
X30067 N30067 N30068 Segment
X30068 N30068 N30069 Segment
X30069 N30069 N30070 Segment
X30070 N30070 N30071 Segment
X30071 N30071 N30072 Segment
X30072 N30072 N30073 Segment
X30073 N30073 N30074 Segment
X30074 N30074 N30075 Segment
X30075 N30075 N30076 Segment
X30076 N30076 N30077 Segment
X30077 N30077 N30078 Segment
X30078 N30078 N30079 Segment
X30079 N30079 N30080 Segment
X30080 N30080 N30081 Segment
X30081 N30081 N30082 Segment
X30082 N30082 N30083 Segment
X30083 N30083 N30084 Segment
X30084 N30084 N30085 Segment
X30085 N30085 N30086 Segment
X30086 N30086 N30087 Segment
X30087 N30087 N30088 Segment
X30088 N30088 N30089 Segment
X30089 N30089 N30090 Segment
X30090 N30090 N30091 Segment
X30091 N30091 N30092 Segment
X30092 N30092 N30093 Segment
X30093 N30093 N30094 Segment
X30094 N30094 N30095 Segment
X30095 N30095 N30096 Segment
X30096 N30096 N30097 Segment
X30097 N30097 N30098 Segment
X30098 N30098 N30099 Segment
X30099 N30099 N30100 Segment
X30100 N30100 N30101 Segment
X30101 N30101 N30102 Segment
X30102 N30102 N30103 Segment
X30103 N30103 N30104 Segment
X30104 N30104 N30105 Segment
X30105 N30105 N30106 Segment
X30106 N30106 N30107 Segment
X30107 N30107 N30108 Segment
X30108 N30108 N30109 Segment
X30109 N30109 N30110 Segment
X30110 N30110 N30111 Segment
X30111 N30111 N30112 Segment
X30112 N30112 N30113 Segment
X30113 N30113 N30114 Segment
X30114 N30114 N30115 Segment
X30115 N30115 N30116 Segment
X30116 N30116 N30117 Segment
X30117 N30117 N30118 Segment
X30118 N30118 N30119 Segment
X30119 N30119 N30120 Segment
X30120 N30120 N30121 Segment
X30121 N30121 N30122 Segment
X30122 N30122 N30123 Segment
X30123 N30123 N30124 Segment
X30124 N30124 N30125 Segment
X30125 N30125 N30126 Segment
X30126 N30126 N30127 Segment
X30127 N30127 N30128 Segment
X30128 N30128 N30129 Segment
X30129 N30129 N30130 Segment
X30130 N30130 N30131 Segment
X30131 N30131 N30132 Segment
X30132 N30132 N30133 Segment
X30133 N30133 N30134 Segment
X30134 N30134 N30135 Segment
X30135 N30135 N30136 Segment
X30136 N30136 N30137 Segment
X30137 N30137 N30138 Segment
X30138 N30138 N30139 Segment
X30139 N30139 N30140 Segment
X30140 N30140 N30141 Segment
X30141 N30141 N30142 Segment
X30142 N30142 N30143 Segment
X30143 N30143 N30144 Segment
X30144 N30144 N30145 Segment
X30145 N30145 N30146 Segment
X30146 N30146 N30147 Segment
X30147 N30147 N30148 Segment
X30148 N30148 N30149 Segment
X30149 N30149 N30150 Segment
X30150 N30150 N30151 Segment
X30151 N30151 N30152 Segment
X30152 N30152 N30153 Segment
X30153 N30153 N30154 Segment
X30154 N30154 N30155 Segment
X30155 N30155 N30156 Segment
X30156 N30156 N30157 Segment
X30157 N30157 N30158 Segment
X30158 N30158 N30159 Segment
X30159 N30159 N30160 Segment
X30160 N30160 N30161 Segment
X30161 N30161 N30162 Segment
X30162 N30162 N30163 Segment
X30163 N30163 N30164 Segment
X30164 N30164 N30165 Segment
X30165 N30165 N30166 Segment
X30166 N30166 N30167 Segment
X30167 N30167 N30168 Segment
X30168 N30168 N30169 Segment
X30169 N30169 N30170 Segment
X30170 N30170 N30171 Segment
X30171 N30171 N30172 Segment
X30172 N30172 N30173 Segment
X30173 N30173 N30174 Segment
X30174 N30174 N30175 Segment
X30175 N30175 N30176 Segment
X30176 N30176 N30177 Segment
X30177 N30177 N30178 Segment
X30178 N30178 N30179 Segment
X30179 N30179 N30180 Segment
X30180 N30180 N30181 Segment
X30181 N30181 N30182 Segment
X30182 N30182 N30183 Segment
X30183 N30183 N30184 Segment
X30184 N30184 N30185 Segment
X30185 N30185 N30186 Segment
X30186 N30186 N30187 Segment
X30187 N30187 N30188 Segment
X30188 N30188 N30189 Segment
X30189 N30189 N30190 Segment
X30190 N30190 N30191 Segment
X30191 N30191 N30192 Segment
X30192 N30192 N30193 Segment
X30193 N30193 N30194 Segment
X30194 N30194 N30195 Segment
X30195 N30195 N30196 Segment
X30196 N30196 N30197 Segment
X30197 N30197 N30198 Segment
X30198 N30198 N30199 Segment
X30199 N30199 N30200 Segment
X30200 N30200 N30201 Segment
X30201 N30201 N30202 Segment
X30202 N30202 N30203 Segment
X30203 N30203 N30204 Segment
X30204 N30204 N30205 Segment
X30205 N30205 N30206 Segment
X30206 N30206 N30207 Segment
X30207 N30207 N30208 Segment
X30208 N30208 N30209 Segment
X30209 N30209 N30210 Segment
X30210 N30210 N30211 Segment
X30211 N30211 N30212 Segment
X30212 N30212 N30213 Segment
X30213 N30213 N30214 Segment
X30214 N30214 N30215 Segment
X30215 N30215 N30216 Segment
X30216 N30216 N30217 Segment
X30217 N30217 N30218 Segment
X30218 N30218 N30219 Segment
X30219 N30219 N30220 Segment
X30220 N30220 N30221 Segment
X30221 N30221 N30222 Segment
X30222 N30222 N30223 Segment
X30223 N30223 N30224 Segment
X30224 N30224 N30225 Segment
X30225 N30225 N30226 Segment
X30226 N30226 N30227 Segment
X30227 N30227 N30228 Segment
X30228 N30228 N30229 Segment
X30229 N30229 N30230 Segment
X30230 N30230 N30231 Segment
X30231 N30231 N30232 Segment
X30232 N30232 N30233 Segment
X30233 N30233 N30234 Segment
X30234 N30234 N30235 Segment
X30235 N30235 N30236 Segment
X30236 N30236 N30237 Segment
X30237 N30237 N30238 Segment
X30238 N30238 N30239 Segment
X30239 N30239 N30240 Segment
X30240 N30240 N30241 Segment
X30241 N30241 N30242 Segment
X30242 N30242 N30243 Segment
X30243 N30243 N30244 Segment
X30244 N30244 N30245 Segment
X30245 N30245 N30246 Segment
X30246 N30246 N30247 Segment
X30247 N30247 N30248 Segment
X30248 N30248 N30249 Segment
X30249 N30249 N30250 Segment
X30250 N30250 N30251 Segment
X30251 N30251 N30252 Segment
X30252 N30252 N30253 Segment
X30253 N30253 N30254 Segment
X30254 N30254 N30255 Segment
X30255 N30255 N30256 Segment
X30256 N30256 N30257 Segment
X30257 N30257 N30258 Segment
X30258 N30258 N30259 Segment
X30259 N30259 N30260 Segment
X30260 N30260 N30261 Segment
X30261 N30261 N30262 Segment
X30262 N30262 N30263 Segment
X30263 N30263 N30264 Segment
X30264 N30264 N30265 Segment
X30265 N30265 N30266 Segment
X30266 N30266 N30267 Segment
X30267 N30267 N30268 Segment
X30268 N30268 N30269 Segment
X30269 N30269 N30270 Segment
X30270 N30270 N30271 Segment
X30271 N30271 N30272 Segment
X30272 N30272 N30273 Segment
X30273 N30273 N30274 Segment
X30274 N30274 N30275 Segment
X30275 N30275 N30276 Segment
X30276 N30276 N30277 Segment
X30277 N30277 N30278 Segment
X30278 N30278 N30279 Segment
X30279 N30279 N30280 Segment
X30280 N30280 N30281 Segment
X30281 N30281 N30282 Segment
X30282 N30282 N30283 Segment
X30283 N30283 N30284 Segment
X30284 N30284 N30285 Segment
X30285 N30285 N30286 Segment
X30286 N30286 N30287 Segment
X30287 N30287 N30288 Segment
X30288 N30288 N30289 Segment
X30289 N30289 N30290 Segment
X30290 N30290 N30291 Segment
X30291 N30291 N30292 Segment
X30292 N30292 N30293 Segment
X30293 N30293 N30294 Segment
X30294 N30294 N30295 Segment
X30295 N30295 N30296 Segment
X30296 N30296 N30297 Segment
X30297 N30297 N30298 Segment
X30298 N30298 N30299 Segment
X30299 N30299 N30300 Segment
X30300 N30300 N30301 Segment
X30301 N30301 N30302 Segment
X30302 N30302 N30303 Segment
X30303 N30303 N30304 Segment
X30304 N30304 N30305 Segment
X30305 N30305 N30306 Segment
X30306 N30306 N30307 Segment
X30307 N30307 N30308 Segment
X30308 N30308 N30309 Segment
X30309 N30309 N30310 Segment
X30310 N30310 N30311 Segment
X30311 N30311 N30312 Segment
X30312 N30312 N30313 Segment
X30313 N30313 N30314 Segment
X30314 N30314 N30315 Segment
X30315 N30315 N30316 Segment
X30316 N30316 N30317 Segment
X30317 N30317 N30318 Segment
X30318 N30318 N30319 Segment
X30319 N30319 N30320 Segment
X30320 N30320 N30321 Segment
X30321 N30321 N30322 Segment
X30322 N30322 N30323 Segment
X30323 N30323 N30324 Segment
X30324 N30324 N30325 Segment
X30325 N30325 N30326 Segment
X30326 N30326 N30327 Segment
X30327 N30327 N30328 Segment
X30328 N30328 N30329 Segment
X30329 N30329 N30330 Segment
X30330 N30330 N30331 Segment
X30331 N30331 N30332 Segment
X30332 N30332 N30333 Segment
X30333 N30333 N30334 Segment
X30334 N30334 N30335 Segment
X30335 N30335 N30336 Segment
X30336 N30336 N30337 Segment
X30337 N30337 N30338 Segment
X30338 N30338 N30339 Segment
X30339 N30339 N30340 Segment
X30340 N30340 N30341 Segment
X30341 N30341 N30342 Segment
X30342 N30342 N30343 Segment
X30343 N30343 N30344 Segment
X30344 N30344 N30345 Segment
X30345 N30345 N30346 Segment
X30346 N30346 N30347 Segment
X30347 N30347 N30348 Segment
X30348 N30348 N30349 Segment
X30349 N30349 N30350 Segment
X30350 N30350 N30351 Segment
X30351 N30351 N30352 Segment
X30352 N30352 N30353 Segment
X30353 N30353 N30354 Segment
X30354 N30354 N30355 Segment
X30355 N30355 N30356 Segment
X30356 N30356 N30357 Segment
X30357 N30357 N30358 Segment
X30358 N30358 N30359 Segment
X30359 N30359 N30360 Segment
X30360 N30360 N30361 Segment
X30361 N30361 N30362 Segment
X30362 N30362 N30363 Segment
X30363 N30363 N30364 Segment
X30364 N30364 N30365 Segment
X30365 N30365 N30366 Segment
X30366 N30366 N30367 Segment
X30367 N30367 N30368 Segment
X30368 N30368 N30369 Segment
X30369 N30369 N30370 Segment
X30370 N30370 N30371 Segment
X30371 N30371 N30372 Segment
X30372 N30372 N30373 Segment
X30373 N30373 N30374 Segment
X30374 N30374 N30375 Segment
X30375 N30375 N30376 Segment
X30376 N30376 N30377 Segment
X30377 N30377 N30378 Segment
X30378 N30378 N30379 Segment
X30379 N30379 N30380 Segment
X30380 N30380 N30381 Segment
X30381 N30381 N30382 Segment
X30382 N30382 N30383 Segment
X30383 N30383 N30384 Segment
X30384 N30384 N30385 Segment
X30385 N30385 N30386 Segment
X30386 N30386 N30387 Segment
X30387 N30387 N30388 Segment
X30388 N30388 N30389 Segment
X30389 N30389 N30390 Segment
X30390 N30390 N30391 Segment
X30391 N30391 N30392 Segment
X30392 N30392 N30393 Segment
X30393 N30393 N30394 Segment
X30394 N30394 N30395 Segment
X30395 N30395 N30396 Segment
X30396 N30396 N30397 Segment
X30397 N30397 N30398 Segment
X30398 N30398 N30399 Segment
X30399 N30399 N30400 Segment
X30400 N30400 N30401 Segment
X30401 N30401 N30402 Segment
X30402 N30402 N30403 Segment
X30403 N30403 N30404 Segment
X30404 N30404 N30405 Segment
X30405 N30405 N30406 Segment
X30406 N30406 N30407 Segment
X30407 N30407 N30408 Segment
X30408 N30408 N30409 Segment
X30409 N30409 N30410 Segment
X30410 N30410 N30411 Segment
X30411 N30411 N30412 Segment
X30412 N30412 N30413 Segment
X30413 N30413 N30414 Segment
X30414 N30414 N30415 Segment
X30415 N30415 N30416 Segment
X30416 N30416 N30417 Segment
X30417 N30417 N30418 Segment
X30418 N30418 N30419 Segment
X30419 N30419 N30420 Segment
X30420 N30420 N30421 Segment
X30421 N30421 N30422 Segment
X30422 N30422 N30423 Segment
X30423 N30423 N30424 Segment
X30424 N30424 N30425 Segment
X30425 N30425 N30426 Segment
X30426 N30426 N30427 Segment
X30427 N30427 N30428 Segment
X30428 N30428 N30429 Segment
X30429 N30429 N30430 Segment
X30430 N30430 N30431 Segment
X30431 N30431 N30432 Segment
X30432 N30432 N30433 Segment
X30433 N30433 N30434 Segment
X30434 N30434 N30435 Segment
X30435 N30435 N30436 Segment
X30436 N30436 N30437 Segment
X30437 N30437 N30438 Segment
X30438 N30438 N30439 Segment
X30439 N30439 N30440 Segment
X30440 N30440 N30441 Segment
X30441 N30441 N30442 Segment
X30442 N30442 N30443 Segment
X30443 N30443 N30444 Segment
X30444 N30444 N30445 Segment
X30445 N30445 N30446 Segment
X30446 N30446 N30447 Segment
X30447 N30447 N30448 Segment
X30448 N30448 N30449 Segment
X30449 N30449 N30450 Segment
X30450 N30450 N30451 Segment
X30451 N30451 N30452 Segment
X30452 N30452 N30453 Segment
X30453 N30453 N30454 Segment
X30454 N30454 N30455 Segment
X30455 N30455 N30456 Segment
X30456 N30456 N30457 Segment
X30457 N30457 N30458 Segment
X30458 N30458 N30459 Segment
X30459 N30459 N30460 Segment
X30460 N30460 N30461 Segment
X30461 N30461 N30462 Segment
X30462 N30462 N30463 Segment
X30463 N30463 N30464 Segment
X30464 N30464 N30465 Segment
X30465 N30465 N30466 Segment
X30466 N30466 N30467 Segment
X30467 N30467 N30468 Segment
X30468 N30468 N30469 Segment
X30469 N30469 N30470 Segment
X30470 N30470 N30471 Segment
X30471 N30471 N30472 Segment
X30472 N30472 N30473 Segment
X30473 N30473 N30474 Segment
X30474 N30474 N30475 Segment
X30475 N30475 N30476 Segment
X30476 N30476 N30477 Segment
X30477 N30477 N30478 Segment
X30478 N30478 N30479 Segment
X30479 N30479 N30480 Segment
X30480 N30480 N30481 Segment
X30481 N30481 N30482 Segment
X30482 N30482 N30483 Segment
X30483 N30483 N30484 Segment
X30484 N30484 N30485 Segment
X30485 N30485 N30486 Segment
X30486 N30486 N30487 Segment
X30487 N30487 N30488 Segment
X30488 N30488 N30489 Segment
X30489 N30489 N30490 Segment
X30490 N30490 N30491 Segment
X30491 N30491 N30492 Segment
X30492 N30492 N30493 Segment
X30493 N30493 N30494 Segment
X30494 N30494 N30495 Segment
X30495 N30495 N30496 Segment
X30496 N30496 N30497 Segment
X30497 N30497 N30498 Segment
X30498 N30498 N30499 Segment
X30499 N30499 N30500 Segment
X30500 N30500 N30501 Segment
X30501 N30501 N30502 Segment
X30502 N30502 N30503 Segment
X30503 N30503 N30504 Segment
X30504 N30504 N30505 Segment
X30505 N30505 N30506 Segment
X30506 N30506 N30507 Segment
X30507 N30507 N30508 Segment
X30508 N30508 N30509 Segment
X30509 N30509 N30510 Segment
X30510 N30510 N30511 Segment
X30511 N30511 N30512 Segment
X30512 N30512 N30513 Segment
X30513 N30513 N30514 Segment
X30514 N30514 N30515 Segment
X30515 N30515 N30516 Segment
X30516 N30516 N30517 Segment
X30517 N30517 N30518 Segment
X30518 N30518 N30519 Segment
X30519 N30519 N30520 Segment
X30520 N30520 N30521 Segment
X30521 N30521 N30522 Segment
X30522 N30522 N30523 Segment
X30523 N30523 N30524 Segment
X30524 N30524 N30525 Segment
X30525 N30525 N30526 Segment
X30526 N30526 N30527 Segment
X30527 N30527 N30528 Segment
X30528 N30528 N30529 Segment
X30529 N30529 N30530 Segment
X30530 N30530 N30531 Segment
X30531 N30531 N30532 Segment
X30532 N30532 N30533 Segment
X30533 N30533 N30534 Segment
X30534 N30534 N30535 Segment
X30535 N30535 N30536 Segment
X30536 N30536 N30537 Segment
X30537 N30537 N30538 Segment
X30538 N30538 N30539 Segment
X30539 N30539 N30540 Segment
X30540 N30540 N30541 Segment
X30541 N30541 N30542 Segment
X30542 N30542 N30543 Segment
X30543 N30543 N30544 Segment
X30544 N30544 N30545 Segment
X30545 N30545 N30546 Segment
X30546 N30546 N30547 Segment
X30547 N30547 N30548 Segment
X30548 N30548 N30549 Segment
X30549 N30549 N30550 Segment
X30550 N30550 N30551 Segment
X30551 N30551 N30552 Segment
X30552 N30552 N30553 Segment
X30553 N30553 N30554 Segment
X30554 N30554 N30555 Segment
X30555 N30555 N30556 Segment
X30556 N30556 N30557 Segment
X30557 N30557 N30558 Segment
X30558 N30558 N30559 Segment
X30559 N30559 N30560 Segment
X30560 N30560 N30561 Segment
X30561 N30561 N30562 Segment
X30562 N30562 N30563 Segment
X30563 N30563 N30564 Segment
X30564 N30564 N30565 Segment
X30565 N30565 N30566 Segment
X30566 N30566 N30567 Segment
X30567 N30567 N30568 Segment
X30568 N30568 N30569 Segment
X30569 N30569 N30570 Segment
X30570 N30570 N30571 Segment
X30571 N30571 N30572 Segment
X30572 N30572 N30573 Segment
X30573 N30573 N30574 Segment
X30574 N30574 N30575 Segment
X30575 N30575 N30576 Segment
X30576 N30576 N30577 Segment
X30577 N30577 N30578 Segment
X30578 N30578 N30579 Segment
X30579 N30579 N30580 Segment
X30580 N30580 N30581 Segment
X30581 N30581 N30582 Segment
X30582 N30582 N30583 Segment
X30583 N30583 N30584 Segment
X30584 N30584 N30585 Segment
X30585 N30585 N30586 Segment
X30586 N30586 N30587 Segment
X30587 N30587 N30588 Segment
X30588 N30588 N30589 Segment
X30589 N30589 N30590 Segment
X30590 N30590 N30591 Segment
X30591 N30591 N30592 Segment
X30592 N30592 N30593 Segment
X30593 N30593 N30594 Segment
X30594 N30594 N30595 Segment
X30595 N30595 N30596 Segment
X30596 N30596 N30597 Segment
X30597 N30597 N30598 Segment
X30598 N30598 N30599 Segment
X30599 N30599 N30600 Segment
X30600 N30600 N30601 Segment
X30601 N30601 N30602 Segment
X30602 N30602 N30603 Segment
X30603 N30603 N30604 Segment
X30604 N30604 N30605 Segment
X30605 N30605 N30606 Segment
X30606 N30606 N30607 Segment
X30607 N30607 N30608 Segment
X30608 N30608 N30609 Segment
X30609 N30609 N30610 Segment
X30610 N30610 N30611 Segment
X30611 N30611 N30612 Segment
X30612 N30612 N30613 Segment
X30613 N30613 N30614 Segment
X30614 N30614 N30615 Segment
X30615 N30615 N30616 Segment
X30616 N30616 N30617 Segment
X30617 N30617 N30618 Segment
X30618 N30618 N30619 Segment
X30619 N30619 N30620 Segment
X30620 N30620 N30621 Segment
X30621 N30621 N30622 Segment
X30622 N30622 N30623 Segment
X30623 N30623 N30624 Segment
X30624 N30624 N30625 Segment
X30625 N30625 N30626 Segment
X30626 N30626 N30627 Segment
X30627 N30627 N30628 Segment
X30628 N30628 N30629 Segment
X30629 N30629 N30630 Segment
X30630 N30630 N30631 Segment
X30631 N30631 N30632 Segment
X30632 N30632 N30633 Segment
X30633 N30633 N30634 Segment
X30634 N30634 N30635 Segment
X30635 N30635 N30636 Segment
X30636 N30636 N30637 Segment
X30637 N30637 N30638 Segment
X30638 N30638 N30639 Segment
X30639 N30639 N30640 Segment
X30640 N30640 N30641 Segment
X30641 N30641 N30642 Segment
X30642 N30642 N30643 Segment
X30643 N30643 N30644 Segment
X30644 N30644 N30645 Segment
X30645 N30645 N30646 Segment
X30646 N30646 N30647 Segment
X30647 N30647 N30648 Segment
X30648 N30648 N30649 Segment
X30649 N30649 N30650 Segment
X30650 N30650 N30651 Segment
X30651 N30651 N30652 Segment
X30652 N30652 N30653 Segment
X30653 N30653 N30654 Segment
X30654 N30654 N30655 Segment
X30655 N30655 N30656 Segment
X30656 N30656 N30657 Segment
X30657 N30657 N30658 Segment
X30658 N30658 N30659 Segment
X30659 N30659 N30660 Segment
X30660 N30660 N30661 Segment
X30661 N30661 N30662 Segment
X30662 N30662 N30663 Segment
X30663 N30663 N30664 Segment
X30664 N30664 N30665 Segment
X30665 N30665 N30666 Segment
X30666 N30666 N30667 Segment
X30667 N30667 N30668 Segment
X30668 N30668 N30669 Segment
X30669 N30669 N30670 Segment
X30670 N30670 N30671 Segment
X30671 N30671 N30672 Segment
X30672 N30672 N30673 Segment
X30673 N30673 N30674 Segment
X30674 N30674 N30675 Segment
X30675 N30675 N30676 Segment
X30676 N30676 N30677 Segment
X30677 N30677 N30678 Segment
X30678 N30678 N30679 Segment
X30679 N30679 N30680 Segment
X30680 N30680 N30681 Segment
X30681 N30681 N30682 Segment
X30682 N30682 N30683 Segment
X30683 N30683 N30684 Segment
X30684 N30684 N30685 Segment
X30685 N30685 N30686 Segment
X30686 N30686 N30687 Segment
X30687 N30687 N30688 Segment
X30688 N30688 N30689 Segment
X30689 N30689 N30690 Segment
X30690 N30690 N30691 Segment
X30691 N30691 N30692 Segment
X30692 N30692 N30693 Segment
X30693 N30693 N30694 Segment
X30694 N30694 N30695 Segment
X30695 N30695 N30696 Segment
X30696 N30696 N30697 Segment
X30697 N30697 N30698 Segment
X30698 N30698 N30699 Segment
X30699 N30699 N30700 Segment
X30700 N30700 N30701 Segment
X30701 N30701 N30702 Segment
X30702 N30702 N30703 Segment
X30703 N30703 N30704 Segment
X30704 N30704 N30705 Segment
X30705 N30705 N30706 Segment
X30706 N30706 N30707 Segment
X30707 N30707 N30708 Segment
X30708 N30708 N30709 Segment
X30709 N30709 N30710 Segment
X30710 N30710 N30711 Segment
X30711 N30711 N30712 Segment
X30712 N30712 N30713 Segment
X30713 N30713 N30714 Segment
X30714 N30714 N30715 Segment
X30715 N30715 N30716 Segment
X30716 N30716 N30717 Segment
X30717 N30717 N30718 Segment
X30718 N30718 N30719 Segment
X30719 N30719 N30720 Segment
X30720 N30720 N30721 Segment
X30721 N30721 N30722 Segment
X30722 N30722 N30723 Segment
X30723 N30723 N30724 Segment
X30724 N30724 N30725 Segment
X30725 N30725 N30726 Segment
X30726 N30726 N30727 Segment
X30727 N30727 N30728 Segment
X30728 N30728 N30729 Segment
X30729 N30729 N30730 Segment
X30730 N30730 N30731 Segment
X30731 N30731 N30732 Segment
X30732 N30732 N30733 Segment
X30733 N30733 N30734 Segment
X30734 N30734 N30735 Segment
X30735 N30735 N30736 Segment
X30736 N30736 N30737 Segment
X30737 N30737 N30738 Segment
X30738 N30738 N30739 Segment
X30739 N30739 N30740 Segment
X30740 N30740 N30741 Segment
X30741 N30741 N30742 Segment
X30742 N30742 N30743 Segment
X30743 N30743 N30744 Segment
X30744 N30744 N30745 Segment
X30745 N30745 N30746 Segment
X30746 N30746 N30747 Segment
X30747 N30747 N30748 Segment
X30748 N30748 N30749 Segment
X30749 N30749 N30750 Segment
X30750 N30750 N30751 Segment
X30751 N30751 N30752 Segment
X30752 N30752 N30753 Segment
X30753 N30753 N30754 Segment
X30754 N30754 N30755 Segment
X30755 N30755 N30756 Segment
X30756 N30756 N30757 Segment
X30757 N30757 N30758 Segment
X30758 N30758 N30759 Segment
X30759 N30759 N30760 Segment
X30760 N30760 N30761 Segment
X30761 N30761 N30762 Segment
X30762 N30762 N30763 Segment
X30763 N30763 N30764 Segment
X30764 N30764 N30765 Segment
X30765 N30765 N30766 Segment
X30766 N30766 N30767 Segment
X30767 N30767 N30768 Segment
X30768 N30768 N30769 Segment
X30769 N30769 N30770 Segment
X30770 N30770 N30771 Segment
X30771 N30771 N30772 Segment
X30772 N30772 N30773 Segment
X30773 N30773 N30774 Segment
X30774 N30774 N30775 Segment
X30775 N30775 N30776 Segment
X30776 N30776 N30777 Segment
X30777 N30777 N30778 Segment
X30778 N30778 N30779 Segment
X30779 N30779 N30780 Segment
X30780 N30780 N30781 Segment
X30781 N30781 N30782 Segment
X30782 N30782 N30783 Segment
X30783 N30783 N30784 Segment
X30784 N30784 N30785 Segment
X30785 N30785 N30786 Segment
X30786 N30786 N30787 Segment
X30787 N30787 N30788 Segment
X30788 N30788 N30789 Segment
X30789 N30789 N30790 Segment
X30790 N30790 N30791 Segment
X30791 N30791 N30792 Segment
X30792 N30792 N30793 Segment
X30793 N30793 N30794 Segment
X30794 N30794 N30795 Segment
X30795 N30795 N30796 Segment
X30796 N30796 N30797 Segment
X30797 N30797 N30798 Segment
X30798 N30798 N30799 Segment
X30799 N30799 N30800 Segment
X30800 N30800 N30801 Segment
X30801 N30801 N30802 Segment
X30802 N30802 N30803 Segment
X30803 N30803 N30804 Segment
X30804 N30804 N30805 Segment
X30805 N30805 N30806 Segment
X30806 N30806 N30807 Segment
X30807 N30807 N30808 Segment
X30808 N30808 N30809 Segment
X30809 N30809 N30810 Segment
X30810 N30810 N30811 Segment
X30811 N30811 N30812 Segment
X30812 N30812 N30813 Segment
X30813 N30813 N30814 Segment
X30814 N30814 N30815 Segment
X30815 N30815 N30816 Segment
X30816 N30816 N30817 Segment
X30817 N30817 N30818 Segment
X30818 N30818 N30819 Segment
X30819 N30819 N30820 Segment
X30820 N30820 N30821 Segment
X30821 N30821 N30822 Segment
X30822 N30822 N30823 Segment
X30823 N30823 N30824 Segment
X30824 N30824 N30825 Segment
X30825 N30825 N30826 Segment
X30826 N30826 N30827 Segment
X30827 N30827 N30828 Segment
X30828 N30828 N30829 Segment
X30829 N30829 N30830 Segment
X30830 N30830 N30831 Segment
X30831 N30831 N30832 Segment
X30832 N30832 N30833 Segment
X30833 N30833 N30834 Segment
X30834 N30834 N30835 Segment
X30835 N30835 N30836 Segment
X30836 N30836 N30837 Segment
X30837 N30837 N30838 Segment
X30838 N30838 N30839 Segment
X30839 N30839 N30840 Segment
X30840 N30840 N30841 Segment
X30841 N30841 N30842 Segment
X30842 N30842 N30843 Segment
X30843 N30843 N30844 Segment
X30844 N30844 N30845 Segment
X30845 N30845 N30846 Segment
X30846 N30846 N30847 Segment
X30847 N30847 N30848 Segment
X30848 N30848 N30849 Segment
X30849 N30849 N30850 Segment
X30850 N30850 N30851 Segment
X30851 N30851 N30852 Segment
X30852 N30852 N30853 Segment
X30853 N30853 N30854 Segment
X30854 N30854 N30855 Segment
X30855 N30855 N30856 Segment
X30856 N30856 N30857 Segment
X30857 N30857 N30858 Segment
X30858 N30858 N30859 Segment
X30859 N30859 N30860 Segment
X30860 N30860 N30861 Segment
X30861 N30861 N30862 Segment
X30862 N30862 N30863 Segment
X30863 N30863 N30864 Segment
X30864 N30864 N30865 Segment
X30865 N30865 N30866 Segment
X30866 N30866 N30867 Segment
X30867 N30867 N30868 Segment
X30868 N30868 N30869 Segment
X30869 N30869 N30870 Segment
X30870 N30870 N30871 Segment
X30871 N30871 N30872 Segment
X30872 N30872 N30873 Segment
X30873 N30873 N30874 Segment
X30874 N30874 N30875 Segment
X30875 N30875 N30876 Segment
X30876 N30876 N30877 Segment
X30877 N30877 N30878 Segment
X30878 N30878 N30879 Segment
X30879 N30879 N30880 Segment
X30880 N30880 N30881 Segment
X30881 N30881 N30882 Segment
X30882 N30882 N30883 Segment
X30883 N30883 N30884 Segment
X30884 N30884 N30885 Segment
X30885 N30885 N30886 Segment
X30886 N30886 N30887 Segment
X30887 N30887 N30888 Segment
X30888 N30888 N30889 Segment
X30889 N30889 N30890 Segment
X30890 N30890 N30891 Segment
X30891 N30891 N30892 Segment
X30892 N30892 N30893 Segment
X30893 N30893 N30894 Segment
X30894 N30894 N30895 Segment
X30895 N30895 N30896 Segment
X30896 N30896 N30897 Segment
X30897 N30897 N30898 Segment
X30898 N30898 N30899 Segment
X30899 N30899 N30900 Segment
X30900 N30900 N30901 Segment
X30901 N30901 N30902 Segment
X30902 N30902 N30903 Segment
X30903 N30903 N30904 Segment
X30904 N30904 N30905 Segment
X30905 N30905 N30906 Segment
X30906 N30906 N30907 Segment
X30907 N30907 N30908 Segment
X30908 N30908 N30909 Segment
X30909 N30909 N30910 Segment
X30910 N30910 N30911 Segment
X30911 N30911 N30912 Segment
X30912 N30912 N30913 Segment
X30913 N30913 N30914 Segment
X30914 N30914 N30915 Segment
X30915 N30915 N30916 Segment
X30916 N30916 N30917 Segment
X30917 N30917 N30918 Segment
X30918 N30918 N30919 Segment
X30919 N30919 N30920 Segment
X30920 N30920 N30921 Segment
X30921 N30921 N30922 Segment
X30922 N30922 N30923 Segment
X30923 N30923 N30924 Segment
X30924 N30924 N30925 Segment
X30925 N30925 N30926 Segment
X30926 N30926 N30927 Segment
X30927 N30927 N30928 Segment
X30928 N30928 N30929 Segment
X30929 N30929 N30930 Segment
X30930 N30930 N30931 Segment
X30931 N30931 N30932 Segment
X30932 N30932 N30933 Segment
X30933 N30933 N30934 Segment
X30934 N30934 N30935 Segment
X30935 N30935 N30936 Segment
X30936 N30936 N30937 Segment
X30937 N30937 N30938 Segment
X30938 N30938 N30939 Segment
X30939 N30939 N30940 Segment
X30940 N30940 N30941 Segment
X30941 N30941 N30942 Segment
X30942 N30942 N30943 Segment
X30943 N30943 N30944 Segment
X30944 N30944 N30945 Segment
X30945 N30945 N30946 Segment
X30946 N30946 N30947 Segment
X30947 N30947 N30948 Segment
X30948 N30948 N30949 Segment
X30949 N30949 N30950 Segment
X30950 N30950 N30951 Segment
X30951 N30951 N30952 Segment
X30952 N30952 N30953 Segment
X30953 N30953 N30954 Segment
X30954 N30954 N30955 Segment
X30955 N30955 N30956 Segment
X30956 N30956 N30957 Segment
X30957 N30957 N30958 Segment
X30958 N30958 N30959 Segment
X30959 N30959 N30960 Segment
X30960 N30960 N30961 Segment
X30961 N30961 N30962 Segment
X30962 N30962 N30963 Segment
X30963 N30963 N30964 Segment
X30964 N30964 N30965 Segment
X30965 N30965 N30966 Segment
X30966 N30966 N30967 Segment
X30967 N30967 N30968 Segment
X30968 N30968 N30969 Segment
X30969 N30969 N30970 Segment
X30970 N30970 N30971 Segment
X30971 N30971 N30972 Segment
X30972 N30972 N30973 Segment
X30973 N30973 N30974 Segment
X30974 N30974 N30975 Segment
X30975 N30975 N30976 Segment
X30976 N30976 N30977 Segment
X30977 N30977 N30978 Segment
X30978 N30978 N30979 Segment
X30979 N30979 N30980 Segment
X30980 N30980 N30981 Segment
X30981 N30981 N30982 Segment
X30982 N30982 N30983 Segment
X30983 N30983 N30984 Segment
X30984 N30984 N30985 Segment
X30985 N30985 N30986 Segment
X30986 N30986 N30987 Segment
X30987 N30987 N30988 Segment
X30988 N30988 N30989 Segment
X30989 N30989 N30990 Segment
X30990 N30990 N30991 Segment
X30991 N30991 N30992 Segment
X30992 N30992 N30993 Segment
X30993 N30993 N30994 Segment
X30994 N30994 N30995 Segment
X30995 N30995 N30996 Segment
X30996 N30996 N30997 Segment
X30997 N30997 N30998 Segment
X30998 N30998 N30999 Segment
X30999 N30999 N31000 Segment
X31000 N31000 N31001 Segment
X31001 N31001 N31002 Segment
X31002 N31002 N31003 Segment
X31003 N31003 N31004 Segment
X31004 N31004 N31005 Segment
X31005 N31005 N31006 Segment
X31006 N31006 N31007 Segment
X31007 N31007 N31008 Segment
X31008 N31008 N31009 Segment
X31009 N31009 N31010 Segment
X31010 N31010 N31011 Segment
X31011 N31011 N31012 Segment
X31012 N31012 N31013 Segment
X31013 N31013 N31014 Segment
X31014 N31014 N31015 Segment
X31015 N31015 N31016 Segment
X31016 N31016 N31017 Segment
X31017 N31017 N31018 Segment
X31018 N31018 N31019 Segment
X31019 N31019 N31020 Segment
X31020 N31020 N31021 Segment
X31021 N31021 N31022 Segment
X31022 N31022 N31023 Segment
X31023 N31023 N31024 Segment
X31024 N31024 N31025 Segment
X31025 N31025 N31026 Segment
X31026 N31026 N31027 Segment
X31027 N31027 N31028 Segment
X31028 N31028 N31029 Segment
X31029 N31029 N31030 Segment
X31030 N31030 N31031 Segment
X31031 N31031 N31032 Segment
X31032 N31032 N31033 Segment
X31033 N31033 N31034 Segment
X31034 N31034 N31035 Segment
X31035 N31035 N31036 Segment
X31036 N31036 N31037 Segment
X31037 N31037 N31038 Segment
X31038 N31038 N31039 Segment
X31039 N31039 N31040 Segment
X31040 N31040 N31041 Segment
X31041 N31041 N31042 Segment
X31042 N31042 N31043 Segment
X31043 N31043 N31044 Segment
X31044 N31044 N31045 Segment
X31045 N31045 N31046 Segment
X31046 N31046 N31047 Segment
X31047 N31047 N31048 Segment
X31048 N31048 N31049 Segment
X31049 N31049 N31050 Segment
X31050 N31050 N31051 Segment
X31051 N31051 N31052 Segment
X31052 N31052 N31053 Segment
X31053 N31053 N31054 Segment
X31054 N31054 N31055 Segment
X31055 N31055 N31056 Segment
X31056 N31056 N31057 Segment
X31057 N31057 N31058 Segment
X31058 N31058 N31059 Segment
X31059 N31059 N31060 Segment
X31060 N31060 N31061 Segment
X31061 N31061 N31062 Segment
X31062 N31062 N31063 Segment
X31063 N31063 N31064 Segment
X31064 N31064 N31065 Segment
X31065 N31065 N31066 Segment
X31066 N31066 N31067 Segment
X31067 N31067 N31068 Segment
X31068 N31068 N31069 Segment
X31069 N31069 N31070 Segment
X31070 N31070 N31071 Segment
X31071 N31071 N31072 Segment
X31072 N31072 N31073 Segment
X31073 N31073 N31074 Segment
X31074 N31074 N31075 Segment
X31075 N31075 N31076 Segment
X31076 N31076 N31077 Segment
X31077 N31077 N31078 Segment
X31078 N31078 N31079 Segment
X31079 N31079 N31080 Segment
X31080 N31080 N31081 Segment
X31081 N31081 N31082 Segment
X31082 N31082 N31083 Segment
X31083 N31083 N31084 Segment
X31084 N31084 N31085 Segment
X31085 N31085 N31086 Segment
X31086 N31086 N31087 Segment
X31087 N31087 N31088 Segment
X31088 N31088 N31089 Segment
X31089 N31089 N31090 Segment
X31090 N31090 N31091 Segment
X31091 N31091 N31092 Segment
X31092 N31092 N31093 Segment
X31093 N31093 N31094 Segment
X31094 N31094 N31095 Segment
X31095 N31095 N31096 Segment
X31096 N31096 N31097 Segment
X31097 N31097 N31098 Segment
X31098 N31098 N31099 Segment
X31099 N31099 N31100 Segment
X31100 N31100 N31101 Segment
X31101 N31101 N31102 Segment
X31102 N31102 N31103 Segment
X31103 N31103 N31104 Segment
X31104 N31104 N31105 Segment
X31105 N31105 N31106 Segment
X31106 N31106 N31107 Segment
X31107 N31107 N31108 Segment
X31108 N31108 N31109 Segment
X31109 N31109 N31110 Segment
X31110 N31110 N31111 Segment
X31111 N31111 N31112 Segment
X31112 N31112 N31113 Segment
X31113 N31113 N31114 Segment
X31114 N31114 N31115 Segment
X31115 N31115 N31116 Segment
X31116 N31116 N31117 Segment
X31117 N31117 N31118 Segment
X31118 N31118 N31119 Segment
X31119 N31119 N31120 Segment
X31120 N31120 N31121 Segment
X31121 N31121 N31122 Segment
X31122 N31122 N31123 Segment
X31123 N31123 N31124 Segment
X31124 N31124 N31125 Segment
X31125 N31125 N31126 Segment
X31126 N31126 N31127 Segment
X31127 N31127 N31128 Segment
X31128 N31128 N31129 Segment
X31129 N31129 N31130 Segment
X31130 N31130 N31131 Segment
X31131 N31131 N31132 Segment
X31132 N31132 N31133 Segment
X31133 N31133 N31134 Segment
X31134 N31134 N31135 Segment
X31135 N31135 N31136 Segment
X31136 N31136 N31137 Segment
X31137 N31137 N31138 Segment
X31138 N31138 N31139 Segment
X31139 N31139 N31140 Segment
X31140 N31140 N31141 Segment
X31141 N31141 N31142 Segment
X31142 N31142 N31143 Segment
X31143 N31143 N31144 Segment
X31144 N31144 N31145 Segment
X31145 N31145 N31146 Segment
X31146 N31146 N31147 Segment
X31147 N31147 N31148 Segment
X31148 N31148 N31149 Segment
X31149 N31149 N31150 Segment
X31150 N31150 N31151 Segment
X31151 N31151 N31152 Segment
X31152 N31152 N31153 Segment
X31153 N31153 N31154 Segment
X31154 N31154 N31155 Segment
X31155 N31155 N31156 Segment
X31156 N31156 N31157 Segment
X31157 N31157 N31158 Segment
X31158 N31158 N31159 Segment
X31159 N31159 N31160 Segment
X31160 N31160 N31161 Segment
X31161 N31161 N31162 Segment
X31162 N31162 N31163 Segment
X31163 N31163 N31164 Segment
X31164 N31164 N31165 Segment
X31165 N31165 N31166 Segment
X31166 N31166 N31167 Segment
X31167 N31167 N31168 Segment
X31168 N31168 N31169 Segment
X31169 N31169 N31170 Segment
X31170 N31170 N31171 Segment
X31171 N31171 N31172 Segment
X31172 N31172 N31173 Segment
X31173 N31173 N31174 Segment
X31174 N31174 N31175 Segment
X31175 N31175 N31176 Segment
X31176 N31176 N31177 Segment
X31177 N31177 N31178 Segment
X31178 N31178 N31179 Segment
X31179 N31179 N31180 Segment
X31180 N31180 N31181 Segment
X31181 N31181 N31182 Segment
X31182 N31182 N31183 Segment
X31183 N31183 N31184 Segment
X31184 N31184 N31185 Segment
X31185 N31185 N31186 Segment
X31186 N31186 N31187 Segment
X31187 N31187 N31188 Segment
X31188 N31188 N31189 Segment
X31189 N31189 N31190 Segment
X31190 N31190 N31191 Segment
X31191 N31191 N31192 Segment
X31192 N31192 N31193 Segment
X31193 N31193 N31194 Segment
X31194 N31194 N31195 Segment
X31195 N31195 N31196 Segment
X31196 N31196 N31197 Segment
X31197 N31197 N31198 Segment
X31198 N31198 N31199 Segment
X31199 N31199 N31200 Segment
X31200 N31200 N31201 Segment
X31201 N31201 N31202 Segment
X31202 N31202 N31203 Segment
X31203 N31203 N31204 Segment
X31204 N31204 N31205 Segment
X31205 N31205 N31206 Segment
X31206 N31206 N31207 Segment
X31207 N31207 N31208 Segment
X31208 N31208 N31209 Segment
X31209 N31209 N31210 Segment
X31210 N31210 N31211 Segment
X31211 N31211 N31212 Segment
X31212 N31212 N31213 Segment
X31213 N31213 N31214 Segment
X31214 N31214 N31215 Segment
X31215 N31215 N31216 Segment
X31216 N31216 N31217 Segment
X31217 N31217 N31218 Segment
X31218 N31218 N31219 Segment
X31219 N31219 N31220 Segment
X31220 N31220 N31221 Segment
X31221 N31221 N31222 Segment
X31222 N31222 N31223 Segment
X31223 N31223 N31224 Segment
X31224 N31224 N31225 Segment
X31225 N31225 N31226 Segment
X31226 N31226 N31227 Segment
X31227 N31227 N31228 Segment
X31228 N31228 N31229 Segment
X31229 N31229 N31230 Segment
X31230 N31230 N31231 Segment
X31231 N31231 N31232 Segment
X31232 N31232 N31233 Segment
X31233 N31233 N31234 Segment
X31234 N31234 N31235 Segment
X31235 N31235 N31236 Segment
X31236 N31236 N31237 Segment
X31237 N31237 N31238 Segment
X31238 N31238 N31239 Segment
X31239 N31239 N31240 Segment
X31240 N31240 N31241 Segment
X31241 N31241 N31242 Segment
X31242 N31242 N31243 Segment
X31243 N31243 N31244 Segment
X31244 N31244 N31245 Segment
X31245 N31245 N31246 Segment
X31246 N31246 N31247 Segment
X31247 N31247 N31248 Segment
X31248 N31248 N31249 Segment
X31249 N31249 N31250 Segment
X31250 N31250 N31251 Segment
X31251 N31251 N31252 Segment
X31252 N31252 N31253 Segment
X31253 N31253 N31254 Segment
X31254 N31254 N31255 Segment
X31255 N31255 N31256 Segment
X31256 N31256 N31257 Segment
X31257 N31257 N31258 Segment
X31258 N31258 N31259 Segment
X31259 N31259 N31260 Segment
X31260 N31260 N31261 Segment
X31261 N31261 N31262 Segment
X31262 N31262 N31263 Segment
X31263 N31263 N31264 Segment
X31264 N31264 N31265 Segment
X31265 N31265 N31266 Segment
X31266 N31266 N31267 Segment
X31267 N31267 N31268 Segment
X31268 N31268 N31269 Segment
X31269 N31269 N31270 Segment
X31270 N31270 N31271 Segment
X31271 N31271 N31272 Segment
X31272 N31272 N31273 Segment
X31273 N31273 N31274 Segment
X31274 N31274 N31275 Segment
X31275 N31275 N31276 Segment
X31276 N31276 N31277 Segment
X31277 N31277 N31278 Segment
X31278 N31278 N31279 Segment
X31279 N31279 N31280 Segment
X31280 N31280 N31281 Segment
X31281 N31281 N31282 Segment
X31282 N31282 N31283 Segment
X31283 N31283 N31284 Segment
X31284 N31284 N31285 Segment
X31285 N31285 N31286 Segment
X31286 N31286 N31287 Segment
X31287 N31287 N31288 Segment
X31288 N31288 N31289 Segment
X31289 N31289 N31290 Segment
X31290 N31290 N31291 Segment
X31291 N31291 N31292 Segment
X31292 N31292 N31293 Segment
X31293 N31293 N31294 Segment
X31294 N31294 N31295 Segment
X31295 N31295 N31296 Segment
X31296 N31296 N31297 Segment
X31297 N31297 N31298 Segment
X31298 N31298 N31299 Segment
X31299 N31299 N31300 Segment
X31300 N31300 N31301 Segment
X31301 N31301 N31302 Segment
X31302 N31302 N31303 Segment
X31303 N31303 N31304 Segment
X31304 N31304 N31305 Segment
X31305 N31305 N31306 Segment
X31306 N31306 N31307 Segment
X31307 N31307 N31308 Segment
X31308 N31308 N31309 Segment
X31309 N31309 N31310 Segment
X31310 N31310 N31311 Segment
X31311 N31311 N31312 Segment
X31312 N31312 N31313 Segment
X31313 N31313 N31314 Segment
X31314 N31314 N31315 Segment
X31315 N31315 N31316 Segment
X31316 N31316 N31317 Segment
X31317 N31317 N31318 Segment
X31318 N31318 N31319 Segment
X31319 N31319 N31320 Segment
X31320 N31320 N31321 Segment
X31321 N31321 N31322 Segment
X31322 N31322 N31323 Segment
X31323 N31323 N31324 Segment
X31324 N31324 N31325 Segment
X31325 N31325 N31326 Segment
X31326 N31326 N31327 Segment
X31327 N31327 N31328 Segment
X31328 N31328 N31329 Segment
X31329 N31329 N31330 Segment
X31330 N31330 N31331 Segment
X31331 N31331 N31332 Segment
X31332 N31332 N31333 Segment
X31333 N31333 N31334 Segment
X31334 N31334 N31335 Segment
X31335 N31335 N31336 Segment
X31336 N31336 N31337 Segment
X31337 N31337 N31338 Segment
X31338 N31338 N31339 Segment
X31339 N31339 N31340 Segment
X31340 N31340 N31341 Segment
X31341 N31341 N31342 Segment
X31342 N31342 N31343 Segment
X31343 N31343 N31344 Segment
X31344 N31344 N31345 Segment
X31345 N31345 N31346 Segment
X31346 N31346 N31347 Segment
X31347 N31347 N31348 Segment
X31348 N31348 N31349 Segment
X31349 N31349 N31350 Segment
X31350 N31350 N31351 Segment
X31351 N31351 N31352 Segment
X31352 N31352 N31353 Segment
X31353 N31353 N31354 Segment
X31354 N31354 N31355 Segment
X31355 N31355 N31356 Segment
X31356 N31356 N31357 Segment
X31357 N31357 N31358 Segment
X31358 N31358 N31359 Segment
X31359 N31359 N31360 Segment
X31360 N31360 N31361 Segment
X31361 N31361 N31362 Segment
X31362 N31362 N31363 Segment
X31363 N31363 N31364 Segment
X31364 N31364 N31365 Segment
X31365 N31365 N31366 Segment
X31366 N31366 N31367 Segment
X31367 N31367 N31368 Segment
X31368 N31368 N31369 Segment
X31369 N31369 N31370 Segment
X31370 N31370 N31371 Segment
X31371 N31371 N31372 Segment
X31372 N31372 N31373 Segment
X31373 N31373 N31374 Segment
X31374 N31374 N31375 Segment
X31375 N31375 N31376 Segment
X31376 N31376 N31377 Segment
X31377 N31377 N31378 Segment
X31378 N31378 N31379 Segment
X31379 N31379 N31380 Segment
X31380 N31380 N31381 Segment
X31381 N31381 N31382 Segment
X31382 N31382 N31383 Segment
X31383 N31383 N31384 Segment
X31384 N31384 N31385 Segment
X31385 N31385 N31386 Segment
X31386 N31386 N31387 Segment
X31387 N31387 N31388 Segment
X31388 N31388 N31389 Segment
X31389 N31389 N31390 Segment
X31390 N31390 N31391 Segment
X31391 N31391 N31392 Segment
X31392 N31392 N31393 Segment
X31393 N31393 N31394 Segment
X31394 N31394 N31395 Segment
X31395 N31395 N31396 Segment
X31396 N31396 N31397 Segment
X31397 N31397 N31398 Segment
X31398 N31398 N31399 Segment
X31399 N31399 N31400 Segment
X31400 N31400 N31401 Segment
X31401 N31401 N31402 Segment
X31402 N31402 N31403 Segment
X31403 N31403 N31404 Segment
X31404 N31404 N31405 Segment
X31405 N31405 N31406 Segment
X31406 N31406 N31407 Segment
X31407 N31407 N31408 Segment
X31408 N31408 N31409 Segment
X31409 N31409 N31410 Segment
X31410 N31410 N31411 Segment
X31411 N31411 N31412 Segment
X31412 N31412 N31413 Segment
X31413 N31413 N31414 Segment
X31414 N31414 N31415 Segment
X31415 N31415 N31416 Segment
X31416 N31416 N31417 Segment
X31417 N31417 N31418 Segment
X31418 N31418 N31419 Segment
X31419 N31419 N31420 Segment
X31420 N31420 N31421 Segment
X31421 N31421 N31422 Segment
X31422 N31422 N31423 Segment
X31423 N31423 N31424 Segment
X31424 N31424 N31425 Segment
X31425 N31425 N31426 Segment
X31426 N31426 N31427 Segment
X31427 N31427 N31428 Segment
X31428 N31428 N31429 Segment
X31429 N31429 N31430 Segment
X31430 N31430 N31431 Segment
X31431 N31431 N31432 Segment
X31432 N31432 N31433 Segment
X31433 N31433 N31434 Segment
X31434 N31434 N31435 Segment
X31435 N31435 N31436 Segment
X31436 N31436 N31437 Segment
X31437 N31437 N31438 Segment
X31438 N31438 N31439 Segment
X31439 N31439 N31440 Segment
X31440 N31440 N31441 Segment
X31441 N31441 N31442 Segment
X31442 N31442 N31443 Segment
X31443 N31443 N31444 Segment
X31444 N31444 N31445 Segment
X31445 N31445 N31446 Segment
X31446 N31446 N31447 Segment
X31447 N31447 N31448 Segment
X31448 N31448 N31449 Segment
X31449 N31449 N31450 Segment
X31450 N31450 N31451 Segment
X31451 N31451 N31452 Segment
X31452 N31452 N31453 Segment
X31453 N31453 N31454 Segment
X31454 N31454 N31455 Segment
X31455 N31455 N31456 Segment
X31456 N31456 N31457 Segment
X31457 N31457 N31458 Segment
X31458 N31458 N31459 Segment
X31459 N31459 N31460 Segment
X31460 N31460 N31461 Segment
X31461 N31461 N31462 Segment
X31462 N31462 N31463 Segment
X31463 N31463 N31464 Segment
X31464 N31464 N31465 Segment
X31465 N31465 N31466 Segment
X31466 N31466 N31467 Segment
X31467 N31467 N31468 Segment
X31468 N31468 N31469 Segment
X31469 N31469 N31470 Segment
X31470 N31470 N31471 Segment
X31471 N31471 N31472 Segment
X31472 N31472 N31473 Segment
X31473 N31473 N31474 Segment
X31474 N31474 N31475 Segment
X31475 N31475 N31476 Segment
X31476 N31476 N31477 Segment
X31477 N31477 N31478 Segment
X31478 N31478 N31479 Segment
X31479 N31479 N31480 Segment
X31480 N31480 N31481 Segment
X31481 N31481 N31482 Segment
X31482 N31482 N31483 Segment
X31483 N31483 N31484 Segment
X31484 N31484 N31485 Segment
X31485 N31485 N31486 Segment
X31486 N31486 N31487 Segment
X31487 N31487 N31488 Segment
X31488 N31488 N31489 Segment
X31489 N31489 N31490 Segment
X31490 N31490 N31491 Segment
X31491 N31491 N31492 Segment
X31492 N31492 N31493 Segment
X31493 N31493 N31494 Segment
X31494 N31494 N31495 Segment
X31495 N31495 N31496 Segment
X31496 N31496 N31497 Segment
X31497 N31497 N31498 Segment
X31498 N31498 N31499 Segment
X31499 N31499 N31500 Segment
X31500 N31500 N31501 Segment
X31501 N31501 N31502 Segment
X31502 N31502 N31503 Segment
X31503 N31503 N31504 Segment
X31504 N31504 N31505 Segment
X31505 N31505 N31506 Segment
X31506 N31506 N31507 Segment
X31507 N31507 N31508 Segment
X31508 N31508 N31509 Segment
X31509 N31509 N31510 Segment
X31510 N31510 N31511 Segment
X31511 N31511 N31512 Segment
X31512 N31512 N31513 Segment
X31513 N31513 N31514 Segment
X31514 N31514 N31515 Segment
X31515 N31515 N31516 Segment
X31516 N31516 N31517 Segment
X31517 N31517 N31518 Segment
X31518 N31518 N31519 Segment
X31519 N31519 N31520 Segment
X31520 N31520 N31521 Segment
X31521 N31521 N31522 Segment
X31522 N31522 N31523 Segment
X31523 N31523 N31524 Segment
X31524 N31524 N31525 Segment
X31525 N31525 N31526 Segment
X31526 N31526 N31527 Segment
X31527 N31527 N31528 Segment
X31528 N31528 N31529 Segment
X31529 N31529 N31530 Segment
X31530 N31530 N31531 Segment
X31531 N31531 N31532 Segment
X31532 N31532 N31533 Segment
X31533 N31533 N31534 Segment
X31534 N31534 N31535 Segment
X31535 N31535 N31536 Segment
X31536 N31536 N31537 Segment
X31537 N31537 N31538 Segment
X31538 N31538 N31539 Segment
X31539 N31539 N31540 Segment
X31540 N31540 N31541 Segment
X31541 N31541 N31542 Segment
X31542 N31542 N31543 Segment
X31543 N31543 N31544 Segment
X31544 N31544 N31545 Segment
X31545 N31545 N31546 Segment
X31546 N31546 N31547 Segment
X31547 N31547 N31548 Segment
X31548 N31548 N31549 Segment
X31549 N31549 N31550 Segment
X31550 N31550 N31551 Segment
X31551 N31551 N31552 Segment
X31552 N31552 N31553 Segment
X31553 N31553 N31554 Segment
X31554 N31554 N31555 Segment
X31555 N31555 N31556 Segment
X31556 N31556 N31557 Segment
X31557 N31557 N31558 Segment
X31558 N31558 N31559 Segment
X31559 N31559 N31560 Segment
X31560 N31560 N31561 Segment
X31561 N31561 N31562 Segment
X31562 N31562 N31563 Segment
X31563 N31563 N31564 Segment
X31564 N31564 N31565 Segment
X31565 N31565 N31566 Segment
X31566 N31566 N31567 Segment
X31567 N31567 N31568 Segment
X31568 N31568 N31569 Segment
X31569 N31569 N31570 Segment
X31570 N31570 N31571 Segment
X31571 N31571 N31572 Segment
X31572 N31572 N31573 Segment
X31573 N31573 N31574 Segment
X31574 N31574 N31575 Segment
X31575 N31575 N31576 Segment
X31576 N31576 N31577 Segment
X31577 N31577 N31578 Segment
X31578 N31578 N31579 Segment
X31579 N31579 N31580 Segment
X31580 N31580 N31581 Segment
X31581 N31581 N31582 Segment
X31582 N31582 N31583 Segment
X31583 N31583 N31584 Segment
X31584 N31584 N31585 Segment
X31585 N31585 N31586 Segment
X31586 N31586 N31587 Segment
X31587 N31587 N31588 Segment
X31588 N31588 N31589 Segment
X31589 N31589 N31590 Segment
X31590 N31590 N31591 Segment
X31591 N31591 N31592 Segment
X31592 N31592 N31593 Segment
X31593 N31593 N31594 Segment
X31594 N31594 N31595 Segment
X31595 N31595 N31596 Segment
X31596 N31596 N31597 Segment
X31597 N31597 N31598 Segment
X31598 N31598 N31599 Segment
X31599 N31599 N31600 Segment
X31600 N31600 N31601 Segment
X31601 N31601 N31602 Segment
X31602 N31602 N31603 Segment
X31603 N31603 N31604 Segment
X31604 N31604 N31605 Segment
X31605 N31605 N31606 Segment
X31606 N31606 N31607 Segment
X31607 N31607 N31608 Segment
X31608 N31608 N31609 Segment
X31609 N31609 N31610 Segment
X31610 N31610 N31611 Segment
X31611 N31611 N31612 Segment
X31612 N31612 N31613 Segment
X31613 N31613 N31614 Segment
X31614 N31614 N31615 Segment
X31615 N31615 N31616 Segment
X31616 N31616 N31617 Segment
X31617 N31617 N31618 Segment
X31618 N31618 N31619 Segment
X31619 N31619 N31620 Segment
X31620 N31620 N31621 Segment
X31621 N31621 N31622 Segment
X31622 N31622 N31623 Segment
X31623 N31623 N31624 Segment
X31624 N31624 N31625 Segment
X31625 N31625 N31626 Segment
X31626 N31626 N31627 Segment
X31627 N31627 N31628 Segment
X31628 N31628 N31629 Segment
X31629 N31629 N31630 Segment
X31630 N31630 N31631 Segment
X31631 N31631 N31632 Segment
X31632 N31632 N31633 Segment
X31633 N31633 N31634 Segment
X31634 N31634 N31635 Segment
X31635 N31635 N31636 Segment
X31636 N31636 N31637 Segment
X31637 N31637 N31638 Segment
X31638 N31638 N31639 Segment
X31639 N31639 N31640 Segment
X31640 N31640 N31641 Segment
X31641 N31641 N31642 Segment
X31642 N31642 N31643 Segment
X31643 N31643 N31644 Segment
X31644 N31644 N31645 Segment
X31645 N31645 N31646 Segment
X31646 N31646 N31647 Segment
X31647 N31647 N31648 Segment
X31648 N31648 N31649 Segment
X31649 N31649 N31650 Segment
X31650 N31650 N31651 Segment
X31651 N31651 N31652 Segment
X31652 N31652 N31653 Segment
X31653 N31653 N31654 Segment
X31654 N31654 N31655 Segment
X31655 N31655 N31656 Segment
X31656 N31656 N31657 Segment
X31657 N31657 N31658 Segment
X31658 N31658 N31659 Segment
X31659 N31659 N31660 Segment
X31660 N31660 N31661 Segment
X31661 N31661 N31662 Segment
X31662 N31662 N31663 Segment
X31663 N31663 N31664 Segment
X31664 N31664 N31665 Segment
X31665 N31665 N31666 Segment
X31666 N31666 N31667 Segment
X31667 N31667 N31668 Segment
X31668 N31668 N31669 Segment
X31669 N31669 N31670 Segment
X31670 N31670 N31671 Segment
X31671 N31671 N31672 Segment
X31672 N31672 N31673 Segment
X31673 N31673 N31674 Segment
X31674 N31674 N31675 Segment
X31675 N31675 N31676 Segment
X31676 N31676 N31677 Segment
X31677 N31677 N31678 Segment
X31678 N31678 N31679 Segment
X31679 N31679 N31680 Segment
X31680 N31680 N31681 Segment
X31681 N31681 N31682 Segment
X31682 N31682 N31683 Segment
X31683 N31683 N31684 Segment
X31684 N31684 N31685 Segment
X31685 N31685 N31686 Segment
X31686 N31686 N31687 Segment
X31687 N31687 N31688 Segment
X31688 N31688 N31689 Segment
X31689 N31689 N31690 Segment
X31690 N31690 N31691 Segment
X31691 N31691 N31692 Segment
X31692 N31692 N31693 Segment
X31693 N31693 N31694 Segment
X31694 N31694 N31695 Segment
X31695 N31695 N31696 Segment
X31696 N31696 N31697 Segment
X31697 N31697 N31698 Segment
X31698 N31698 N31699 Segment
X31699 N31699 N31700 Segment
X31700 N31700 N31701 Segment
X31701 N31701 N31702 Segment
X31702 N31702 N31703 Segment
X31703 N31703 N31704 Segment
X31704 N31704 N31705 Segment
X31705 N31705 N31706 Segment
X31706 N31706 N31707 Segment
X31707 N31707 N31708 Segment
X31708 N31708 N31709 Segment
X31709 N31709 N31710 Segment
X31710 N31710 N31711 Segment
X31711 N31711 N31712 Segment
X31712 N31712 N31713 Segment
X31713 N31713 N31714 Segment
X31714 N31714 N31715 Segment
X31715 N31715 N31716 Segment
X31716 N31716 N31717 Segment
X31717 N31717 N31718 Segment
X31718 N31718 N31719 Segment
X31719 N31719 N31720 Segment
X31720 N31720 N31721 Segment
X31721 N31721 N31722 Segment
X31722 N31722 N31723 Segment
X31723 N31723 N31724 Segment
X31724 N31724 N31725 Segment
X31725 N31725 N31726 Segment
X31726 N31726 N31727 Segment
X31727 N31727 N31728 Segment
X31728 N31728 N31729 Segment
X31729 N31729 N31730 Segment
X31730 N31730 N31731 Segment
X31731 N31731 N31732 Segment
X31732 N31732 N31733 Segment
X31733 N31733 N31734 Segment
X31734 N31734 N31735 Segment
X31735 N31735 N31736 Segment
X31736 N31736 N31737 Segment
X31737 N31737 N31738 Segment
X31738 N31738 N31739 Segment
X31739 N31739 N31740 Segment
X31740 N31740 N31741 Segment
X31741 N31741 N31742 Segment
X31742 N31742 N31743 Segment
X31743 N31743 N31744 Segment
X31744 N31744 N31745 Segment
X31745 N31745 N31746 Segment
X31746 N31746 N31747 Segment
X31747 N31747 N31748 Segment
X31748 N31748 N31749 Segment
X31749 N31749 N31750 Segment
X31750 N31750 N31751 Segment
X31751 N31751 N31752 Segment
X31752 N31752 N31753 Segment
X31753 N31753 N31754 Segment
X31754 N31754 N31755 Segment
X31755 N31755 N31756 Segment
X31756 N31756 N31757 Segment
X31757 N31757 N31758 Segment
X31758 N31758 N31759 Segment
X31759 N31759 N31760 Segment
X31760 N31760 N31761 Segment
X31761 N31761 N31762 Segment
X31762 N31762 N31763 Segment
X31763 N31763 N31764 Segment
X31764 N31764 N31765 Segment
X31765 N31765 N31766 Segment
X31766 N31766 N31767 Segment
X31767 N31767 N31768 Segment
X31768 N31768 N31769 Segment
X31769 N31769 N31770 Segment
X31770 N31770 N31771 Segment
X31771 N31771 N31772 Segment
X31772 N31772 N31773 Segment
X31773 N31773 N31774 Segment
X31774 N31774 N31775 Segment
X31775 N31775 N31776 Segment
X31776 N31776 N31777 Segment
X31777 N31777 N31778 Segment
X31778 N31778 N31779 Segment
X31779 N31779 N31780 Segment
X31780 N31780 N31781 Segment
X31781 N31781 N31782 Segment
X31782 N31782 N31783 Segment
X31783 N31783 N31784 Segment
X31784 N31784 N31785 Segment
X31785 N31785 N31786 Segment
X31786 N31786 N31787 Segment
X31787 N31787 N31788 Segment
X31788 N31788 N31789 Segment
X31789 N31789 N31790 Segment
X31790 N31790 N31791 Segment
X31791 N31791 N31792 Segment
X31792 N31792 N31793 Segment
X31793 N31793 N31794 Segment
X31794 N31794 N31795 Segment
X31795 N31795 N31796 Segment
X31796 N31796 N31797 Segment
X31797 N31797 N31798 Segment
X31798 N31798 N31799 Segment
X31799 N31799 N31800 Segment
X31800 N31800 N31801 Segment
X31801 N31801 N31802 Segment
X31802 N31802 N31803 Segment
X31803 N31803 N31804 Segment
X31804 N31804 N31805 Segment
X31805 N31805 N31806 Segment
X31806 N31806 N31807 Segment
X31807 N31807 N31808 Segment
X31808 N31808 N31809 Segment
X31809 N31809 N31810 Segment
X31810 N31810 N31811 Segment
X31811 N31811 N31812 Segment
X31812 N31812 N31813 Segment
X31813 N31813 N31814 Segment
X31814 N31814 N31815 Segment
X31815 N31815 N31816 Segment
X31816 N31816 N31817 Segment
X31817 N31817 N31818 Segment
X31818 N31818 N31819 Segment
X31819 N31819 N31820 Segment
X31820 N31820 N31821 Segment
X31821 N31821 N31822 Segment
X31822 N31822 N31823 Segment
X31823 N31823 N31824 Segment
X31824 N31824 N31825 Segment
X31825 N31825 N31826 Segment
X31826 N31826 N31827 Segment
X31827 N31827 N31828 Segment
X31828 N31828 N31829 Segment
X31829 N31829 N31830 Segment
X31830 N31830 N31831 Segment
X31831 N31831 N31832 Segment
X31832 N31832 N31833 Segment
X31833 N31833 N31834 Segment
X31834 N31834 N31835 Segment
X31835 N31835 N31836 Segment
X31836 N31836 N31837 Segment
X31837 N31837 N31838 Segment
X31838 N31838 N31839 Segment
X31839 N31839 N31840 Segment
X31840 N31840 N31841 Segment
X31841 N31841 N31842 Segment
X31842 N31842 N31843 Segment
X31843 N31843 N31844 Segment
X31844 N31844 N31845 Segment
X31845 N31845 N31846 Segment
X31846 N31846 N31847 Segment
X31847 N31847 N31848 Segment
X31848 N31848 N31849 Segment
X31849 N31849 N31850 Segment
X31850 N31850 N31851 Segment
X31851 N31851 N31852 Segment
X31852 N31852 N31853 Segment
X31853 N31853 N31854 Segment
X31854 N31854 N31855 Segment
X31855 N31855 N31856 Segment
X31856 N31856 N31857 Segment
X31857 N31857 N31858 Segment
X31858 N31858 N31859 Segment
X31859 N31859 N31860 Segment
X31860 N31860 N31861 Segment
X31861 N31861 N31862 Segment
X31862 N31862 N31863 Segment
X31863 N31863 N31864 Segment
X31864 N31864 N31865 Segment
X31865 N31865 N31866 Segment
X31866 N31866 N31867 Segment
X31867 N31867 N31868 Segment
X31868 N31868 N31869 Segment
X31869 N31869 N31870 Segment
X31870 N31870 N31871 Segment
X31871 N31871 N31872 Segment
X31872 N31872 N31873 Segment
X31873 N31873 N31874 Segment
X31874 N31874 N31875 Segment
X31875 N31875 N31876 Segment
X31876 N31876 N31877 Segment
X31877 N31877 N31878 Segment
X31878 N31878 N31879 Segment
X31879 N31879 N31880 Segment
X31880 N31880 N31881 Segment
X31881 N31881 N31882 Segment
X31882 N31882 N31883 Segment
X31883 N31883 N31884 Segment
X31884 N31884 N31885 Segment
X31885 N31885 N31886 Segment
X31886 N31886 N31887 Segment
X31887 N31887 N31888 Segment
X31888 N31888 N31889 Segment
X31889 N31889 N31890 Segment
X31890 N31890 N31891 Segment
X31891 N31891 N31892 Segment
X31892 N31892 N31893 Segment
X31893 N31893 N31894 Segment
X31894 N31894 N31895 Segment
X31895 N31895 N31896 Segment
X31896 N31896 N31897 Segment
X31897 N31897 N31898 Segment
X31898 N31898 N31899 Segment
X31899 N31899 N31900 Segment
X31900 N31900 N31901 Segment
X31901 N31901 N31902 Segment
X31902 N31902 N31903 Segment
X31903 N31903 N31904 Segment
X31904 N31904 N31905 Segment
X31905 N31905 N31906 Segment
X31906 N31906 N31907 Segment
X31907 N31907 N31908 Segment
X31908 N31908 N31909 Segment
X31909 N31909 N31910 Segment
X31910 N31910 N31911 Segment
X31911 N31911 N31912 Segment
X31912 N31912 N31913 Segment
X31913 N31913 N31914 Segment
X31914 N31914 N31915 Segment
X31915 N31915 N31916 Segment
X31916 N31916 N31917 Segment
X31917 N31917 N31918 Segment
X31918 N31918 N31919 Segment
X31919 N31919 N31920 Segment
X31920 N31920 N31921 Segment
X31921 N31921 N31922 Segment
X31922 N31922 N31923 Segment
X31923 N31923 N31924 Segment
X31924 N31924 N31925 Segment
X31925 N31925 N31926 Segment
X31926 N31926 N31927 Segment
X31927 N31927 N31928 Segment
X31928 N31928 N31929 Segment
X31929 N31929 N31930 Segment
X31930 N31930 N31931 Segment
X31931 N31931 N31932 Segment
X31932 N31932 N31933 Segment
X31933 N31933 N31934 Segment
X31934 N31934 N31935 Segment
X31935 N31935 N31936 Segment
X31936 N31936 N31937 Segment
X31937 N31937 N31938 Segment
X31938 N31938 N31939 Segment
X31939 N31939 N31940 Segment
X31940 N31940 N31941 Segment
X31941 N31941 N31942 Segment
X31942 N31942 N31943 Segment
X31943 N31943 N31944 Segment
X31944 N31944 N31945 Segment
X31945 N31945 N31946 Segment
X31946 N31946 N31947 Segment
X31947 N31947 N31948 Segment
X31948 N31948 N31949 Segment
X31949 N31949 N31950 Segment
X31950 N31950 N31951 Segment
X31951 N31951 N31952 Segment
X31952 N31952 N31953 Segment
X31953 N31953 N31954 Segment
X31954 N31954 N31955 Segment
X31955 N31955 N31956 Segment
X31956 N31956 N31957 Segment
X31957 N31957 N31958 Segment
X31958 N31958 N31959 Segment
X31959 N31959 N31960 Segment
X31960 N31960 N31961 Segment
X31961 N31961 N31962 Segment
X31962 N31962 N31963 Segment
X31963 N31963 N31964 Segment
X31964 N31964 N31965 Segment
X31965 N31965 N31966 Segment
X31966 N31966 N31967 Segment
X31967 N31967 N31968 Segment
X31968 N31968 N31969 Segment
X31969 N31969 N31970 Segment
X31970 N31970 N31971 Segment
X31971 N31971 N31972 Segment
X31972 N31972 N31973 Segment
X31973 N31973 N31974 Segment
X31974 N31974 N31975 Segment
X31975 N31975 N31976 Segment
X31976 N31976 N31977 Segment
X31977 N31977 N31978 Segment
X31978 N31978 N31979 Segment
X31979 N31979 N31980 Segment
X31980 N31980 N31981 Segment
X31981 N31981 N31982 Segment
X31982 N31982 N31983 Segment
X31983 N31983 N31984 Segment
X31984 N31984 N31985 Segment
X31985 N31985 N31986 Segment
X31986 N31986 N31987 Segment
X31987 N31987 N31988 Segment
X31988 N31988 N31989 Segment
X31989 N31989 N31990 Segment
X31990 N31990 N31991 Segment
X31991 N31991 N31992 Segment
X31992 N31992 N31993 Segment
X31993 N31993 N31994 Segment
X31994 N31994 N31995 Segment
X31995 N31995 N31996 Segment
X31996 N31996 N31997 Segment
X31997 N31997 N31998 Segment
X31998 N31998 N31999 Segment
X31999 N31999 N32000 Segment
X32000 N32000 N32001 Segment
X32001 N32001 N32002 Segment
X32002 N32002 N32003 Segment
X32003 N32003 N32004 Segment
X32004 N32004 N32005 Segment
X32005 N32005 N32006 Segment
X32006 N32006 N32007 Segment
X32007 N32007 N32008 Segment
X32008 N32008 N32009 Segment
X32009 N32009 N32010 Segment
X32010 N32010 N32011 Segment
X32011 N32011 N32012 Segment
X32012 N32012 N32013 Segment
X32013 N32013 N32014 Segment
X32014 N32014 N32015 Segment
X32015 N32015 N32016 Segment
X32016 N32016 N32017 Segment
X32017 N32017 N32018 Segment
X32018 N32018 N32019 Segment
X32019 N32019 N32020 Segment
X32020 N32020 N32021 Segment
X32021 N32021 N32022 Segment
X32022 N32022 N32023 Segment
X32023 N32023 N32024 Segment
X32024 N32024 N32025 Segment
X32025 N32025 N32026 Segment
X32026 N32026 N32027 Segment
X32027 N32027 N32028 Segment
X32028 N32028 N32029 Segment
X32029 N32029 N32030 Segment
X32030 N32030 N32031 Segment
X32031 N32031 N32032 Segment
X32032 N32032 N32033 Segment
X32033 N32033 N32034 Segment
X32034 N32034 N32035 Segment
X32035 N32035 N32036 Segment
X32036 N32036 N32037 Segment
X32037 N32037 N32038 Segment
X32038 N32038 N32039 Segment
X32039 N32039 N32040 Segment
X32040 N32040 N32041 Segment
X32041 N32041 N32042 Segment
X32042 N32042 N32043 Segment
X32043 N32043 N32044 Segment
X32044 N32044 N32045 Segment
X32045 N32045 N32046 Segment
X32046 N32046 N32047 Segment
X32047 N32047 N32048 Segment
X32048 N32048 N32049 Segment
X32049 N32049 N32050 Segment
X32050 N32050 N32051 Segment
X32051 N32051 N32052 Segment
X32052 N32052 N32053 Segment
X32053 N32053 N32054 Segment
X32054 N32054 N32055 Segment
X32055 N32055 N32056 Segment
X32056 N32056 N32057 Segment
X32057 N32057 N32058 Segment
X32058 N32058 N32059 Segment
X32059 N32059 N32060 Segment
X32060 N32060 N32061 Segment
X32061 N32061 N32062 Segment
X32062 N32062 N32063 Segment
X32063 N32063 N32064 Segment
X32064 N32064 N32065 Segment
X32065 N32065 N32066 Segment
X32066 N32066 N32067 Segment
X32067 N32067 N32068 Segment
X32068 N32068 N32069 Segment
X32069 N32069 N32070 Segment
X32070 N32070 N32071 Segment
X32071 N32071 N32072 Segment
X32072 N32072 N32073 Segment
X32073 N32073 N32074 Segment
X32074 N32074 N32075 Segment
X32075 N32075 N32076 Segment
X32076 N32076 N32077 Segment
X32077 N32077 N32078 Segment
X32078 N32078 N32079 Segment
X32079 N32079 N32080 Segment
X32080 N32080 N32081 Segment
X32081 N32081 N32082 Segment
X32082 N32082 N32083 Segment
X32083 N32083 N32084 Segment
X32084 N32084 N32085 Segment
X32085 N32085 N32086 Segment
X32086 N32086 N32087 Segment
X32087 N32087 N32088 Segment
X32088 N32088 N32089 Segment
X32089 N32089 N32090 Segment
X32090 N32090 N32091 Segment
X32091 N32091 N32092 Segment
X32092 N32092 N32093 Segment
X32093 N32093 N32094 Segment
X32094 N32094 N32095 Segment
X32095 N32095 N32096 Segment
X32096 N32096 N32097 Segment
X32097 N32097 N32098 Segment
X32098 N32098 N32099 Segment
X32099 N32099 N32100 Segment
X32100 N32100 N32101 Segment
X32101 N32101 N32102 Segment
X32102 N32102 N32103 Segment
X32103 N32103 N32104 Segment
X32104 N32104 N32105 Segment
X32105 N32105 N32106 Segment
X32106 N32106 N32107 Segment
X32107 N32107 N32108 Segment
X32108 N32108 N32109 Segment
X32109 N32109 N32110 Segment
X32110 N32110 N32111 Segment
X32111 N32111 N32112 Segment
X32112 N32112 N32113 Segment
X32113 N32113 N32114 Segment
X32114 N32114 N32115 Segment
X32115 N32115 N32116 Segment
X32116 N32116 N32117 Segment
X32117 N32117 N32118 Segment
X32118 N32118 N32119 Segment
X32119 N32119 N32120 Segment
X32120 N32120 N32121 Segment
X32121 N32121 N32122 Segment
X32122 N32122 N32123 Segment
X32123 N32123 N32124 Segment
X32124 N32124 N32125 Segment
X32125 N32125 N32126 Segment
X32126 N32126 N32127 Segment
X32127 N32127 N32128 Segment
X32128 N32128 N32129 Segment
X32129 N32129 N32130 Segment
X32130 N32130 N32131 Segment
X32131 N32131 N32132 Segment
X32132 N32132 N32133 Segment
X32133 N32133 N32134 Segment
X32134 N32134 N32135 Segment
X32135 N32135 N32136 Segment
X32136 N32136 N32137 Segment
X32137 N32137 N32138 Segment
X32138 N32138 N32139 Segment
X32139 N32139 N32140 Segment
X32140 N32140 N32141 Segment
X32141 N32141 N32142 Segment
X32142 N32142 N32143 Segment
X32143 N32143 N32144 Segment
X32144 N32144 N32145 Segment
X32145 N32145 N32146 Segment
X32146 N32146 N32147 Segment
X32147 N32147 N32148 Segment
X32148 N32148 N32149 Segment
X32149 N32149 N32150 Segment
X32150 N32150 N32151 Segment
X32151 N32151 N32152 Segment
X32152 N32152 N32153 Segment
X32153 N32153 N32154 Segment
X32154 N32154 N32155 Segment
X32155 N32155 N32156 Segment
X32156 N32156 N32157 Segment
X32157 N32157 N32158 Segment
X32158 N32158 N32159 Segment
X32159 N32159 N32160 Segment
X32160 N32160 N32161 Segment
X32161 N32161 N32162 Segment
X32162 N32162 N32163 Segment
X32163 N32163 N32164 Segment
X32164 N32164 N32165 Segment
X32165 N32165 N32166 Segment
X32166 N32166 N32167 Segment
X32167 N32167 N32168 Segment
X32168 N32168 N32169 Segment
X32169 N32169 N32170 Segment
X32170 N32170 N32171 Segment
X32171 N32171 N32172 Segment
X32172 N32172 N32173 Segment
X32173 N32173 N32174 Segment
X32174 N32174 N32175 Segment
X32175 N32175 N32176 Segment
X32176 N32176 N32177 Segment
X32177 N32177 N32178 Segment
X32178 N32178 N32179 Segment
X32179 N32179 N32180 Segment
X32180 N32180 N32181 Segment
X32181 N32181 N32182 Segment
X32182 N32182 N32183 Segment
X32183 N32183 N32184 Segment
X32184 N32184 N32185 Segment
X32185 N32185 N32186 Segment
X32186 N32186 N32187 Segment
X32187 N32187 N32188 Segment
X32188 N32188 N32189 Segment
X32189 N32189 N32190 Segment
X32190 N32190 N32191 Segment
X32191 N32191 N32192 Segment
X32192 N32192 N32193 Segment
X32193 N32193 N32194 Segment
X32194 N32194 N32195 Segment
X32195 N32195 N32196 Segment
X32196 N32196 N32197 Segment
X32197 N32197 N32198 Segment
X32198 N32198 N32199 Segment
X32199 N32199 N32200 Segment
X32200 N32200 N32201 Segment
X32201 N32201 N32202 Segment
X32202 N32202 N32203 Segment
X32203 N32203 N32204 Segment
X32204 N32204 N32205 Segment
X32205 N32205 N32206 Segment
X32206 N32206 N32207 Segment
X32207 N32207 N32208 Segment
X32208 N32208 N32209 Segment
X32209 N32209 N32210 Segment
X32210 N32210 N32211 Segment
X32211 N32211 N32212 Segment
X32212 N32212 N32213 Segment
X32213 N32213 N32214 Segment
X32214 N32214 N32215 Segment
X32215 N32215 N32216 Segment
X32216 N32216 N32217 Segment
X32217 N32217 N32218 Segment
X32218 N32218 N32219 Segment
X32219 N32219 N32220 Segment
X32220 N32220 N32221 Segment
X32221 N32221 N32222 Segment
X32222 N32222 N32223 Segment
X32223 N32223 N32224 Segment
X32224 N32224 N32225 Segment
X32225 N32225 N32226 Segment
X32226 N32226 N32227 Segment
X32227 N32227 N32228 Segment
X32228 N32228 N32229 Segment
X32229 N32229 N32230 Segment
X32230 N32230 N32231 Segment
X32231 N32231 N32232 Segment
X32232 N32232 N32233 Segment
X32233 N32233 N32234 Segment
X32234 N32234 N32235 Segment
X32235 N32235 N32236 Segment
X32236 N32236 N32237 Segment
X32237 N32237 N32238 Segment
X32238 N32238 N32239 Segment
X32239 N32239 N32240 Segment
X32240 N32240 N32241 Segment
X32241 N32241 N32242 Segment
X32242 N32242 N32243 Segment
X32243 N32243 N32244 Segment
X32244 N32244 N32245 Segment
X32245 N32245 N32246 Segment
X32246 N32246 N32247 Segment
X32247 N32247 N32248 Segment
X32248 N32248 N32249 Segment
X32249 N32249 N32250 Segment
X32250 N32250 N32251 Segment
X32251 N32251 N32252 Segment
X32252 N32252 N32253 Segment
X32253 N32253 N32254 Segment
X32254 N32254 N32255 Segment
X32255 N32255 N32256 Segment
X32256 N32256 N32257 Segment
X32257 N32257 N32258 Segment
X32258 N32258 N32259 Segment
X32259 N32259 N32260 Segment
X32260 N32260 N32261 Segment
X32261 N32261 N32262 Segment
X32262 N32262 N32263 Segment
X32263 N32263 N32264 Segment
X32264 N32264 N32265 Segment
X32265 N32265 N32266 Segment
X32266 N32266 N32267 Segment
X32267 N32267 N32268 Segment
X32268 N32268 N32269 Segment
X32269 N32269 N32270 Segment
X32270 N32270 N32271 Segment
X32271 N32271 N32272 Segment
X32272 N32272 N32273 Segment
X32273 N32273 N32274 Segment
X32274 N32274 N32275 Segment
X32275 N32275 N32276 Segment
X32276 N32276 N32277 Segment
X32277 N32277 N32278 Segment
X32278 N32278 N32279 Segment
X32279 N32279 N32280 Segment
X32280 N32280 N32281 Segment
X32281 N32281 N32282 Segment
X32282 N32282 N32283 Segment
X32283 N32283 N32284 Segment
X32284 N32284 N32285 Segment
X32285 N32285 N32286 Segment
X32286 N32286 N32287 Segment
X32287 N32287 N32288 Segment
X32288 N32288 N32289 Segment
X32289 N32289 N32290 Segment
X32290 N32290 N32291 Segment
X32291 N32291 N32292 Segment
X32292 N32292 N32293 Segment
X32293 N32293 N32294 Segment
X32294 N32294 N32295 Segment
X32295 N32295 N32296 Segment
X32296 N32296 N32297 Segment
X32297 N32297 N32298 Segment
X32298 N32298 N32299 Segment
X32299 N32299 N32300 Segment
X32300 N32300 N32301 Segment
X32301 N32301 N32302 Segment
X32302 N32302 N32303 Segment
X32303 N32303 N32304 Segment
X32304 N32304 N32305 Segment
X32305 N32305 N32306 Segment
X32306 N32306 N32307 Segment
X32307 N32307 N32308 Segment
X32308 N32308 N32309 Segment
X32309 N32309 N32310 Segment
X32310 N32310 N32311 Segment
X32311 N32311 N32312 Segment
X32312 N32312 N32313 Segment
X32313 N32313 N32314 Segment
X32314 N32314 N32315 Segment
X32315 N32315 N32316 Segment
X32316 N32316 N32317 Segment
X32317 N32317 N32318 Segment
X32318 N32318 N32319 Segment
X32319 N32319 N32320 Segment
X32320 N32320 N32321 Segment
X32321 N32321 N32322 Segment
X32322 N32322 N32323 Segment
X32323 N32323 N32324 Segment
X32324 N32324 N32325 Segment
X32325 N32325 N32326 Segment
X32326 N32326 N32327 Segment
X32327 N32327 N32328 Segment
X32328 N32328 N32329 Segment
X32329 N32329 N32330 Segment
X32330 N32330 N32331 Segment
X32331 N32331 N32332 Segment
X32332 N32332 N32333 Segment
X32333 N32333 N32334 Segment
X32334 N32334 N32335 Segment
X32335 N32335 N32336 Segment
X32336 N32336 N32337 Segment
X32337 N32337 N32338 Segment
X32338 N32338 N32339 Segment
X32339 N32339 N32340 Segment
X32340 N32340 N32341 Segment
X32341 N32341 N32342 Segment
X32342 N32342 N32343 Segment
X32343 N32343 N32344 Segment
X32344 N32344 N32345 Segment
X32345 N32345 N32346 Segment
X32346 N32346 N32347 Segment
X32347 N32347 N32348 Segment
X32348 N32348 N32349 Segment
X32349 N32349 N32350 Segment
X32350 N32350 N32351 Segment
X32351 N32351 N32352 Segment
X32352 N32352 N32353 Segment
X32353 N32353 N32354 Segment
X32354 N32354 N32355 Segment
X32355 N32355 N32356 Segment
X32356 N32356 N32357 Segment
X32357 N32357 N32358 Segment
X32358 N32358 N32359 Segment
X32359 N32359 N32360 Segment
X32360 N32360 N32361 Segment
X32361 N32361 N32362 Segment
X32362 N32362 N32363 Segment
X32363 N32363 N32364 Segment
X32364 N32364 N32365 Segment
X32365 N32365 N32366 Segment
X32366 N32366 N32367 Segment
X32367 N32367 N32368 Segment
X32368 N32368 N32369 Segment
X32369 N32369 N32370 Segment
X32370 N32370 N32371 Segment
X32371 N32371 N32372 Segment
X32372 N32372 N32373 Segment
X32373 N32373 N32374 Segment
X32374 N32374 N32375 Segment
X32375 N32375 N32376 Segment
X32376 N32376 N32377 Segment
X32377 N32377 N32378 Segment
X32378 N32378 N32379 Segment
X32379 N32379 N32380 Segment
X32380 N32380 N32381 Segment
X32381 N32381 N32382 Segment
X32382 N32382 N32383 Segment
X32383 N32383 N32384 Segment
X32384 N32384 N32385 Segment
X32385 N32385 N32386 Segment
X32386 N32386 N32387 Segment
X32387 N32387 N32388 Segment
X32388 N32388 N32389 Segment
X32389 N32389 N32390 Segment
X32390 N32390 N32391 Segment
X32391 N32391 N32392 Segment
X32392 N32392 N32393 Segment
X32393 N32393 N32394 Segment
X32394 N32394 N32395 Segment
X32395 N32395 N32396 Segment
X32396 N32396 N32397 Segment
X32397 N32397 N32398 Segment
X32398 N32398 N32399 Segment
X32399 N32399 N32400 Segment
X32400 N32400 N32401 Segment
X32401 N32401 N32402 Segment
X32402 N32402 N32403 Segment
X32403 N32403 N32404 Segment
X32404 N32404 N32405 Segment
X32405 N32405 N32406 Segment
X32406 N32406 N32407 Segment
X32407 N32407 N32408 Segment
X32408 N32408 N32409 Segment
X32409 N32409 N32410 Segment
X32410 N32410 N32411 Segment
X32411 N32411 N32412 Segment
X32412 N32412 N32413 Segment
X32413 N32413 N32414 Segment
X32414 N32414 N32415 Segment
X32415 N32415 N32416 Segment
X32416 N32416 N32417 Segment
X32417 N32417 N32418 Segment
X32418 N32418 N32419 Segment
X32419 N32419 N32420 Segment
X32420 N32420 N32421 Segment
X32421 N32421 N32422 Segment
X32422 N32422 N32423 Segment
X32423 N32423 N32424 Segment
X32424 N32424 N32425 Segment
X32425 N32425 N32426 Segment
X32426 N32426 N32427 Segment
X32427 N32427 N32428 Segment
X32428 N32428 N32429 Segment
X32429 N32429 N32430 Segment
X32430 N32430 N32431 Segment
X32431 N32431 N32432 Segment
X32432 N32432 N32433 Segment
X32433 N32433 N32434 Segment
X32434 N32434 N32435 Segment
X32435 N32435 N32436 Segment
X32436 N32436 N32437 Segment
X32437 N32437 N32438 Segment
X32438 N32438 N32439 Segment
X32439 N32439 N32440 Segment
X32440 N32440 N32441 Segment
X32441 N32441 N32442 Segment
X32442 N32442 N32443 Segment
X32443 N32443 N32444 Segment
X32444 N32444 N32445 Segment
X32445 N32445 N32446 Segment
X32446 N32446 N32447 Segment
X32447 N32447 N32448 Segment
X32448 N32448 N32449 Segment
X32449 N32449 N32450 Segment
X32450 N32450 N32451 Segment
X32451 N32451 N32452 Segment
X32452 N32452 N32453 Segment
X32453 N32453 N32454 Segment
X32454 N32454 N32455 Segment
X32455 N32455 N32456 Segment
X32456 N32456 N32457 Segment
X32457 N32457 N32458 Segment
X32458 N32458 N32459 Segment
X32459 N32459 N32460 Segment
X32460 N32460 N32461 Segment
X32461 N32461 N32462 Segment
X32462 N32462 N32463 Segment
X32463 N32463 N32464 Segment
X32464 N32464 N32465 Segment
X32465 N32465 N32466 Segment
X32466 N32466 N32467 Segment
X32467 N32467 N32468 Segment
X32468 N32468 N32469 Segment
X32469 N32469 N32470 Segment
X32470 N32470 N32471 Segment
X32471 N32471 N32472 Segment
X32472 N32472 N32473 Segment
X32473 N32473 N32474 Segment
X32474 N32474 N32475 Segment
X32475 N32475 N32476 Segment
X32476 N32476 N32477 Segment
X32477 N32477 N32478 Segment
X32478 N32478 N32479 Segment
X32479 N32479 N32480 Segment
X32480 N32480 N32481 Segment
X32481 N32481 N32482 Segment
X32482 N32482 N32483 Segment
X32483 N32483 N32484 Segment
X32484 N32484 N32485 Segment
X32485 N32485 N32486 Segment
X32486 N32486 N32487 Segment
X32487 N32487 N32488 Segment
X32488 N32488 N32489 Segment
X32489 N32489 N32490 Segment
X32490 N32490 N32491 Segment
X32491 N32491 N32492 Segment
X32492 N32492 N32493 Segment
X32493 N32493 N32494 Segment
X32494 N32494 N32495 Segment
X32495 N32495 N32496 Segment
X32496 N32496 N32497 Segment
X32497 N32497 N32498 Segment
X32498 N32498 N32499 Segment
X32499 N32499 N32500 Segment
X32500 N32500 N32501 Segment
X32501 N32501 N32502 Segment
X32502 N32502 N32503 Segment
X32503 N32503 N32504 Segment
X32504 N32504 N32505 Segment
X32505 N32505 N32506 Segment
X32506 N32506 N32507 Segment
X32507 N32507 N32508 Segment
X32508 N32508 N32509 Segment
X32509 N32509 N32510 Segment
X32510 N32510 N32511 Segment
X32511 N32511 N32512 Segment
X32512 N32512 N32513 Segment
X32513 N32513 N32514 Segment
X32514 N32514 N32515 Segment
X32515 N32515 N32516 Segment
X32516 N32516 N32517 Segment
X32517 N32517 N32518 Segment
X32518 N32518 N32519 Segment
X32519 N32519 N32520 Segment
X32520 N32520 N32521 Segment
X32521 N32521 N32522 Segment
X32522 N32522 N32523 Segment
X32523 N32523 N32524 Segment
X32524 N32524 N32525 Segment
X32525 N32525 N32526 Segment
X32526 N32526 N32527 Segment
X32527 N32527 N32528 Segment
X32528 N32528 N32529 Segment
X32529 N32529 N32530 Segment
X32530 N32530 N32531 Segment
X32531 N32531 N32532 Segment
X32532 N32532 N32533 Segment
X32533 N32533 N32534 Segment
X32534 N32534 N32535 Segment
X32535 N32535 N32536 Segment
X32536 N32536 N32537 Segment
X32537 N32537 N32538 Segment
X32538 N32538 N32539 Segment
X32539 N32539 N32540 Segment
X32540 N32540 N32541 Segment
X32541 N32541 N32542 Segment
X32542 N32542 N32543 Segment
X32543 N32543 N32544 Segment
X32544 N32544 N32545 Segment
X32545 N32545 N32546 Segment
X32546 N32546 N32547 Segment
X32547 N32547 N32548 Segment
X32548 N32548 N32549 Segment
X32549 N32549 N32550 Segment
X32550 N32550 N32551 Segment
X32551 N32551 N32552 Segment
X32552 N32552 N32553 Segment
X32553 N32553 N32554 Segment
X32554 N32554 N32555 Segment
X32555 N32555 N32556 Segment
X32556 N32556 N32557 Segment
X32557 N32557 N32558 Segment
X32558 N32558 N32559 Segment
X32559 N32559 N32560 Segment
X32560 N32560 N32561 Segment
X32561 N32561 N32562 Segment
X32562 N32562 N32563 Segment
X32563 N32563 N32564 Segment
X32564 N32564 N32565 Segment
X32565 N32565 N32566 Segment
X32566 N32566 N32567 Segment
X32567 N32567 N32568 Segment
X32568 N32568 N32569 Segment
X32569 N32569 N32570 Segment
X32570 N32570 N32571 Segment
X32571 N32571 N32572 Segment
X32572 N32572 N32573 Segment
X32573 N32573 N32574 Segment
X32574 N32574 N32575 Segment
X32575 N32575 N32576 Segment
X32576 N32576 N32577 Segment
X32577 N32577 N32578 Segment
X32578 N32578 N32579 Segment
X32579 N32579 N32580 Segment
X32580 N32580 N32581 Segment
X32581 N32581 N32582 Segment
X32582 N32582 N32583 Segment
X32583 N32583 N32584 Segment
X32584 N32584 N32585 Segment
X32585 N32585 N32586 Segment
X32586 N32586 N32587 Segment
X32587 N32587 N32588 Segment
X32588 N32588 N32589 Segment
X32589 N32589 N32590 Segment
X32590 N32590 N32591 Segment
X32591 N32591 N32592 Segment
X32592 N32592 N32593 Segment
X32593 N32593 N32594 Segment
X32594 N32594 N32595 Segment
X32595 N32595 N32596 Segment
X32596 N32596 N32597 Segment
X32597 N32597 N32598 Segment
X32598 N32598 N32599 Segment
X32599 N32599 N32600 Segment
X32600 N32600 N32601 Segment
X32601 N32601 N32602 Segment
X32602 N32602 N32603 Segment
X32603 N32603 N32604 Segment
X32604 N32604 N32605 Segment
X32605 N32605 N32606 Segment
X32606 N32606 N32607 Segment
X32607 N32607 N32608 Segment
X32608 N32608 N32609 Segment
X32609 N32609 N32610 Segment
X32610 N32610 N32611 Segment
X32611 N32611 N32612 Segment
X32612 N32612 N32613 Segment
X32613 N32613 N32614 Segment
X32614 N32614 N32615 Segment
X32615 N32615 N32616 Segment
X32616 N32616 N32617 Segment
X32617 N32617 N32618 Segment
X32618 N32618 N32619 Segment
X32619 N32619 N32620 Segment
X32620 N32620 N32621 Segment
X32621 N32621 N32622 Segment
X32622 N32622 N32623 Segment
X32623 N32623 N32624 Segment
X32624 N32624 N32625 Segment
X32625 N32625 N32626 Segment
X32626 N32626 N32627 Segment
X32627 N32627 N32628 Segment
X32628 N32628 N32629 Segment
X32629 N32629 N32630 Segment
X32630 N32630 N32631 Segment
X32631 N32631 N32632 Segment
X32632 N32632 N32633 Segment
X32633 N32633 N32634 Segment
X32634 N32634 N32635 Segment
X32635 N32635 N32636 Segment
X32636 N32636 N32637 Segment
X32637 N32637 N32638 Segment
X32638 N32638 N32639 Segment
X32639 N32639 N32640 Segment
X32640 N32640 N32641 Segment
X32641 N32641 N32642 Segment
X32642 N32642 N32643 Segment
X32643 N32643 N32644 Segment
X32644 N32644 N32645 Segment
X32645 N32645 N32646 Segment
X32646 N32646 N32647 Segment
X32647 N32647 N32648 Segment
X32648 N32648 N32649 Segment
X32649 N32649 N32650 Segment
X32650 N32650 N32651 Segment
X32651 N32651 N32652 Segment
X32652 N32652 N32653 Segment
X32653 N32653 N32654 Segment
X32654 N32654 N32655 Segment
X32655 N32655 N32656 Segment
X32656 N32656 N32657 Segment
X32657 N32657 N32658 Segment
X32658 N32658 N32659 Segment
X32659 N32659 N32660 Segment
X32660 N32660 N32661 Segment
X32661 N32661 N32662 Segment
X32662 N32662 N32663 Segment
X32663 N32663 N32664 Segment
X32664 N32664 N32665 Segment
X32665 N32665 N32666 Segment
X32666 N32666 N32667 Segment
X32667 N32667 N32668 Segment
X32668 N32668 N32669 Segment
X32669 N32669 N32670 Segment
X32670 N32670 N32671 Segment
X32671 N32671 N32672 Segment
X32672 N32672 N32673 Segment
X32673 N32673 N32674 Segment
X32674 N32674 N32675 Segment
X32675 N32675 N32676 Segment
X32676 N32676 N32677 Segment
X32677 N32677 N32678 Segment
X32678 N32678 N32679 Segment
X32679 N32679 N32680 Segment
X32680 N32680 N32681 Segment
X32681 N32681 N32682 Segment
X32682 N32682 N32683 Segment
X32683 N32683 N32684 Segment
X32684 N32684 N32685 Segment
X32685 N32685 N32686 Segment
X32686 N32686 N32687 Segment
X32687 N32687 N32688 Segment
X32688 N32688 N32689 Segment
X32689 N32689 N32690 Segment
X32690 N32690 N32691 Segment
X32691 N32691 N32692 Segment
X32692 N32692 N32693 Segment
X32693 N32693 N32694 Segment
X32694 N32694 N32695 Segment
X32695 N32695 N32696 Segment
X32696 N32696 N32697 Segment
X32697 N32697 N32698 Segment
X32698 N32698 N32699 Segment
X32699 N32699 N32700 Segment
X32700 N32700 N32701 Segment
X32701 N32701 N32702 Segment
X32702 N32702 N32703 Segment
X32703 N32703 N32704 Segment
X32704 N32704 N32705 Segment
X32705 N32705 N32706 Segment
X32706 N32706 N32707 Segment
X32707 N32707 N32708 Segment
X32708 N32708 N32709 Segment
X32709 N32709 N32710 Segment
X32710 N32710 N32711 Segment
X32711 N32711 N32712 Segment
X32712 N32712 N32713 Segment
X32713 N32713 N32714 Segment
X32714 N32714 N32715 Segment
X32715 N32715 N32716 Segment
X32716 N32716 N32717 Segment
X32717 N32717 N32718 Segment
X32718 N32718 N32719 Segment
X32719 N32719 N32720 Segment
X32720 N32720 N32721 Segment
X32721 N32721 N32722 Segment
X32722 N32722 N32723 Segment
X32723 N32723 N32724 Segment
X32724 N32724 N32725 Segment
X32725 N32725 N32726 Segment
X32726 N32726 N32727 Segment
X32727 N32727 N32728 Segment
X32728 N32728 N32729 Segment
X32729 N32729 N32730 Segment
X32730 N32730 N32731 Segment
X32731 N32731 N32732 Segment
X32732 N32732 N32733 Segment
X32733 N32733 N32734 Segment
X32734 N32734 N32735 Segment
X32735 N32735 N32736 Segment
X32736 N32736 N32737 Segment
X32737 N32737 N32738 Segment
X32738 N32738 N32739 Segment
X32739 N32739 N32740 Segment
X32740 N32740 N32741 Segment
X32741 N32741 N32742 Segment
X32742 N32742 N32743 Segment
X32743 N32743 N32744 Segment
X32744 N32744 N32745 Segment
X32745 N32745 N32746 Segment
X32746 N32746 N32747 Segment
X32747 N32747 N32748 Segment
X32748 N32748 N32749 Segment
X32749 N32749 N32750 Segment
X32750 N32750 N32751 Segment
X32751 N32751 N32752 Segment
X32752 N32752 N32753 Segment
X32753 N32753 N32754 Segment
X32754 N32754 N32755 Segment
X32755 N32755 N32756 Segment
X32756 N32756 N32757 Segment
X32757 N32757 N32758 Segment
X32758 N32758 N32759 Segment
X32759 N32759 N32760 Segment
X32760 N32760 N32761 Segment
X32761 N32761 N32762 Segment
X32762 N32762 N32763 Segment
X32763 N32763 N32764 Segment
X32764 N32764 N32765 Segment
X32765 N32765 N32766 Segment
X32766 N32766 N32767 Segment
X32767 N32767 N32768 Segment
X32768 N32768 N32769 Segment
X32769 N32769 N32770 Segment
X32770 N32770 N32771 Segment
X32771 N32771 N32772 Segment
X32772 N32772 N32773 Segment
X32773 N32773 N32774 Segment
X32774 N32774 N32775 Segment
X32775 N32775 N32776 Segment
X32776 N32776 N32777 Segment
X32777 N32777 N32778 Segment
X32778 N32778 N32779 Segment
X32779 N32779 N32780 Segment
X32780 N32780 N32781 Segment
X32781 N32781 N32782 Segment
X32782 N32782 N32783 Segment
X32783 N32783 N32784 Segment
X32784 N32784 N32785 Segment
X32785 N32785 N32786 Segment
X32786 N32786 N32787 Segment
X32787 N32787 N32788 Segment
X32788 N32788 N32789 Segment
X32789 N32789 N32790 Segment
X32790 N32790 N32791 Segment
X32791 N32791 N32792 Segment
X32792 N32792 N32793 Segment
X32793 N32793 N32794 Segment
X32794 N32794 N32795 Segment
X32795 N32795 N32796 Segment
X32796 N32796 N32797 Segment
X32797 N32797 N32798 Segment
X32798 N32798 N32799 Segment
X32799 N32799 N32800 Segment
X32800 N32800 N32801 Segment
X32801 N32801 N32802 Segment
X32802 N32802 N32803 Segment
X32803 N32803 N32804 Segment
X32804 N32804 N32805 Segment
X32805 N32805 N32806 Segment
X32806 N32806 N32807 Segment
X32807 N32807 N32808 Segment
X32808 N32808 N32809 Segment
X32809 N32809 N32810 Segment
X32810 N32810 N32811 Segment
X32811 N32811 N32812 Segment
X32812 N32812 N32813 Segment
X32813 N32813 N32814 Segment
X32814 N32814 N32815 Segment
X32815 N32815 N32816 Segment
X32816 N32816 N32817 Segment
X32817 N32817 N32818 Segment
X32818 N32818 N32819 Segment
X32819 N32819 N32820 Segment
X32820 N32820 N32821 Segment
X32821 N32821 N32822 Segment
X32822 N32822 N32823 Segment
X32823 N32823 N32824 Segment
X32824 N32824 N32825 Segment
X32825 N32825 N32826 Segment
X32826 N32826 N32827 Segment
X32827 N32827 N32828 Segment
X32828 N32828 N32829 Segment
X32829 N32829 N32830 Segment
X32830 N32830 N32831 Segment
X32831 N32831 N32832 Segment
X32832 N32832 N32833 Segment
X32833 N32833 N32834 Segment
X32834 N32834 N32835 Segment
X32835 N32835 N32836 Segment
X32836 N32836 N32837 Segment
X32837 N32837 N32838 Segment
X32838 N32838 N32839 Segment
X32839 N32839 N32840 Segment
X32840 N32840 N32841 Segment
X32841 N32841 N32842 Segment
X32842 N32842 N32843 Segment
X32843 N32843 N32844 Segment
X32844 N32844 N32845 Segment
X32845 N32845 N32846 Segment
X32846 N32846 N32847 Segment
X32847 N32847 N32848 Segment
X32848 N32848 N32849 Segment
X32849 N32849 N32850 Segment
X32850 N32850 N32851 Segment
X32851 N32851 N32852 Segment
X32852 N32852 N32853 Segment
X32853 N32853 N32854 Segment
X32854 N32854 N32855 Segment
X32855 N32855 N32856 Segment
X32856 N32856 N32857 Segment
X32857 N32857 N32858 Segment
X32858 N32858 N32859 Segment
X32859 N32859 N32860 Segment
X32860 N32860 N32861 Segment
X32861 N32861 N32862 Segment
X32862 N32862 N32863 Segment
X32863 N32863 N32864 Segment
X32864 N32864 N32865 Segment
X32865 N32865 N32866 Segment
X32866 N32866 N32867 Segment
X32867 N32867 N32868 Segment
X32868 N32868 N32869 Segment
X32869 N32869 N32870 Segment
X32870 N32870 N32871 Segment
X32871 N32871 N32872 Segment
X32872 N32872 N32873 Segment
X32873 N32873 N32874 Segment
X32874 N32874 N32875 Segment
X32875 N32875 N32876 Segment
X32876 N32876 N32877 Segment
X32877 N32877 N32878 Segment
X32878 N32878 N32879 Segment
X32879 N32879 N32880 Segment
X32880 N32880 N32881 Segment
X32881 N32881 N32882 Segment
X32882 N32882 N32883 Segment
X32883 N32883 N32884 Segment
X32884 N32884 N32885 Segment
X32885 N32885 N32886 Segment
X32886 N32886 N32887 Segment
X32887 N32887 N32888 Segment
X32888 N32888 N32889 Segment
X32889 N32889 N32890 Segment
X32890 N32890 N32891 Segment
X32891 N32891 N32892 Segment
X32892 N32892 N32893 Segment
X32893 N32893 N32894 Segment
X32894 N32894 N32895 Segment
X32895 N32895 N32896 Segment
X32896 N32896 N32897 Segment
X32897 N32897 N32898 Segment
X32898 N32898 N32899 Segment
X32899 N32899 N32900 Segment
X32900 N32900 N32901 Segment
X32901 N32901 N32902 Segment
X32902 N32902 N32903 Segment
X32903 N32903 N32904 Segment
X32904 N32904 N32905 Segment
X32905 N32905 N32906 Segment
X32906 N32906 N32907 Segment
X32907 N32907 N32908 Segment
X32908 N32908 N32909 Segment
X32909 N32909 N32910 Segment
X32910 N32910 N32911 Segment
X32911 N32911 N32912 Segment
X32912 N32912 N32913 Segment
X32913 N32913 N32914 Segment
X32914 N32914 N32915 Segment
X32915 N32915 N32916 Segment
X32916 N32916 N32917 Segment
X32917 N32917 N32918 Segment
X32918 N32918 N32919 Segment
X32919 N32919 N32920 Segment
X32920 N32920 N32921 Segment
X32921 N32921 N32922 Segment
X32922 N32922 N32923 Segment
X32923 N32923 N32924 Segment
X32924 N32924 N32925 Segment
X32925 N32925 N32926 Segment
X32926 N32926 N32927 Segment
X32927 N32927 N32928 Segment
X32928 N32928 N32929 Segment
X32929 N32929 N32930 Segment
X32930 N32930 N32931 Segment
X32931 N32931 N32932 Segment
X32932 N32932 N32933 Segment
X32933 N32933 N32934 Segment
X32934 N32934 N32935 Segment
X32935 N32935 N32936 Segment
X32936 N32936 N32937 Segment
X32937 N32937 N32938 Segment
X32938 N32938 N32939 Segment
X32939 N32939 N32940 Segment
X32940 N32940 N32941 Segment
X32941 N32941 N32942 Segment
X32942 N32942 N32943 Segment
X32943 N32943 N32944 Segment
X32944 N32944 N32945 Segment
X32945 N32945 N32946 Segment
X32946 N32946 N32947 Segment
X32947 N32947 N32948 Segment
X32948 N32948 N32949 Segment
X32949 N32949 N32950 Segment
X32950 N32950 N32951 Segment
X32951 N32951 N32952 Segment
X32952 N32952 N32953 Segment
X32953 N32953 N32954 Segment
X32954 N32954 N32955 Segment
X32955 N32955 N32956 Segment
X32956 N32956 N32957 Segment
X32957 N32957 N32958 Segment
X32958 N32958 N32959 Segment
X32959 N32959 N32960 Segment
X32960 N32960 N32961 Segment
X32961 N32961 N32962 Segment
X32962 N32962 N32963 Segment
X32963 N32963 N32964 Segment
X32964 N32964 N32965 Segment
X32965 N32965 N32966 Segment
X32966 N32966 N32967 Segment
X32967 N32967 N32968 Segment
X32968 N32968 N32969 Segment
X32969 N32969 N32970 Segment
X32970 N32970 N32971 Segment
X32971 N32971 N32972 Segment
X32972 N32972 N32973 Segment
X32973 N32973 N32974 Segment
X32974 N32974 N32975 Segment
X32975 N32975 N32976 Segment
X32976 N32976 N32977 Segment
X32977 N32977 N32978 Segment
X32978 N32978 N32979 Segment
X32979 N32979 N32980 Segment
X32980 N32980 N32981 Segment
X32981 N32981 N32982 Segment
X32982 N32982 N32983 Segment
X32983 N32983 N32984 Segment
X32984 N32984 N32985 Segment
X32985 N32985 N32986 Segment
X32986 N32986 N32987 Segment
X32987 N32987 N32988 Segment
X32988 N32988 N32989 Segment
X32989 N32989 N32990 Segment
X32990 N32990 N32991 Segment
X32991 N32991 N32992 Segment
X32992 N32992 N32993 Segment
X32993 N32993 N32994 Segment
X32994 N32994 N32995 Segment
X32995 N32995 N32996 Segment
X32996 N32996 N32997 Segment
X32997 N32997 N32998 Segment
X32998 N32998 N32999 Segment
X32999 N32999 N33000 Segment
X33000 N33000 N33001 Segment
X33001 N33001 N33002 Segment
X33002 N33002 N33003 Segment
X33003 N33003 N33004 Segment
X33004 N33004 N33005 Segment
X33005 N33005 N33006 Segment
X33006 N33006 N33007 Segment
X33007 N33007 N33008 Segment
X33008 N33008 N33009 Segment
X33009 N33009 N33010 Segment
X33010 N33010 N33011 Segment
X33011 N33011 N33012 Segment
X33012 N33012 N33013 Segment
X33013 N33013 N33014 Segment
X33014 N33014 N33015 Segment
X33015 N33015 N33016 Segment
X33016 N33016 N33017 Segment
X33017 N33017 N33018 Segment
X33018 N33018 N33019 Segment
X33019 N33019 N33020 Segment
X33020 N33020 N33021 Segment
X33021 N33021 N33022 Segment
X33022 N33022 N33023 Segment
X33023 N33023 N33024 Segment
X33024 N33024 N33025 Segment
X33025 N33025 N33026 Segment
X33026 N33026 N33027 Segment
X33027 N33027 N33028 Segment
X33028 N33028 N33029 Segment
X33029 N33029 N33030 Segment
X33030 N33030 N33031 Segment
X33031 N33031 N33032 Segment
X33032 N33032 N33033 Segment
X33033 N33033 N33034 Segment
X33034 N33034 N33035 Segment
X33035 N33035 N33036 Segment
X33036 N33036 N33037 Segment
X33037 N33037 N33038 Segment
X33038 N33038 N33039 Segment
X33039 N33039 N33040 Segment
X33040 N33040 N33041 Segment
X33041 N33041 N33042 Segment
X33042 N33042 N33043 Segment
X33043 N33043 N33044 Segment
X33044 N33044 N33045 Segment
X33045 N33045 N33046 Segment
X33046 N33046 N33047 Segment
X33047 N33047 N33048 Segment
X33048 N33048 N33049 Segment
X33049 N33049 N33050 Segment
X33050 N33050 N33051 Segment
X33051 N33051 N33052 Segment
X33052 N33052 N33053 Segment
X33053 N33053 N33054 Segment
X33054 N33054 N33055 Segment
X33055 N33055 N33056 Segment
X33056 N33056 N33057 Segment
X33057 N33057 N33058 Segment
X33058 N33058 N33059 Segment
X33059 N33059 N33060 Segment
X33060 N33060 N33061 Segment
X33061 N33061 N33062 Segment
X33062 N33062 N33063 Segment
X33063 N33063 N33064 Segment
X33064 N33064 N33065 Segment
X33065 N33065 N33066 Segment
X33066 N33066 N33067 Segment
X33067 N33067 N33068 Segment
X33068 N33068 N33069 Segment
X33069 N33069 N33070 Segment
X33070 N33070 N33071 Segment
X33071 N33071 N33072 Segment
X33072 N33072 N33073 Segment
X33073 N33073 N33074 Segment
X33074 N33074 N33075 Segment
X33075 N33075 N33076 Segment
X33076 N33076 N33077 Segment
X33077 N33077 N33078 Segment
X33078 N33078 N33079 Segment
X33079 N33079 N33080 Segment
X33080 N33080 N33081 Segment
X33081 N33081 N33082 Segment
X33082 N33082 N33083 Segment
X33083 N33083 N33084 Segment
X33084 N33084 N33085 Segment
X33085 N33085 N33086 Segment
X33086 N33086 N33087 Segment
X33087 N33087 N33088 Segment
X33088 N33088 N33089 Segment
X33089 N33089 N33090 Segment
X33090 N33090 N33091 Segment
X33091 N33091 N33092 Segment
X33092 N33092 N33093 Segment
X33093 N33093 N33094 Segment
X33094 N33094 N33095 Segment
X33095 N33095 N33096 Segment
X33096 N33096 N33097 Segment
X33097 N33097 N33098 Segment
X33098 N33098 N33099 Segment
X33099 N33099 N33100 Segment
X33100 N33100 N33101 Segment
X33101 N33101 N33102 Segment
X33102 N33102 N33103 Segment
X33103 N33103 N33104 Segment
X33104 N33104 N33105 Segment
X33105 N33105 N33106 Segment
X33106 N33106 N33107 Segment
X33107 N33107 N33108 Segment
X33108 N33108 N33109 Segment
X33109 N33109 N33110 Segment
X33110 N33110 N33111 Segment
X33111 N33111 N33112 Segment
X33112 N33112 N33113 Segment
X33113 N33113 N33114 Segment
X33114 N33114 N33115 Segment
X33115 N33115 N33116 Segment
X33116 N33116 N33117 Segment
X33117 N33117 N33118 Segment
X33118 N33118 N33119 Segment
X33119 N33119 N33120 Segment
X33120 N33120 N33121 Segment
X33121 N33121 N33122 Segment
X33122 N33122 N33123 Segment
X33123 N33123 N33124 Segment
X33124 N33124 N33125 Segment
X33125 N33125 N33126 Segment
X33126 N33126 N33127 Segment
X33127 N33127 N33128 Segment
X33128 N33128 N33129 Segment
X33129 N33129 N33130 Segment
X33130 N33130 N33131 Segment
X33131 N33131 N33132 Segment
X33132 N33132 N33133 Segment
X33133 N33133 N33134 Segment
X33134 N33134 N33135 Segment
X33135 N33135 N33136 Segment
X33136 N33136 N33137 Segment
X33137 N33137 N33138 Segment
X33138 N33138 N33139 Segment
X33139 N33139 N33140 Segment
X33140 N33140 N33141 Segment
X33141 N33141 N33142 Segment
X33142 N33142 N33143 Segment
X33143 N33143 N33144 Segment
X33144 N33144 N33145 Segment
X33145 N33145 N33146 Segment
X33146 N33146 N33147 Segment
X33147 N33147 N33148 Segment
X33148 N33148 N33149 Segment
X33149 N33149 N33150 Segment
X33150 N33150 N33151 Segment
X33151 N33151 N33152 Segment
X33152 N33152 N33153 Segment
X33153 N33153 N33154 Segment
X33154 N33154 N33155 Segment
X33155 N33155 N33156 Segment
X33156 N33156 N33157 Segment
X33157 N33157 N33158 Segment
X33158 N33158 N33159 Segment
X33159 N33159 N33160 Segment
X33160 N33160 N33161 Segment
X33161 N33161 N33162 Segment
X33162 N33162 N33163 Segment
X33163 N33163 N33164 Segment
X33164 N33164 N33165 Segment
X33165 N33165 N33166 Segment
X33166 N33166 N33167 Segment
X33167 N33167 N33168 Segment
X33168 N33168 N33169 Segment
X33169 N33169 N33170 Segment
X33170 N33170 N33171 Segment
X33171 N33171 N33172 Segment
X33172 N33172 N33173 Segment
X33173 N33173 N33174 Segment
X33174 N33174 N33175 Segment
X33175 N33175 N33176 Segment
X33176 N33176 N33177 Segment
X33177 N33177 N33178 Segment
X33178 N33178 N33179 Segment
X33179 N33179 N33180 Segment
X33180 N33180 N33181 Segment
X33181 N33181 N33182 Segment
X33182 N33182 N33183 Segment
X33183 N33183 N33184 Segment
X33184 N33184 N33185 Segment
X33185 N33185 N33186 Segment
X33186 N33186 N33187 Segment
X33187 N33187 N33188 Segment
X33188 N33188 N33189 Segment
X33189 N33189 N33190 Segment
X33190 N33190 N33191 Segment
X33191 N33191 N33192 Segment
X33192 N33192 N33193 Segment
X33193 N33193 N33194 Segment
X33194 N33194 N33195 Segment
X33195 N33195 N33196 Segment
X33196 N33196 N33197 Segment
X33197 N33197 N33198 Segment
X33198 N33198 N33199 Segment
X33199 N33199 N33200 Segment
X33200 N33200 N33201 Segment
X33201 N33201 N33202 Segment
X33202 N33202 N33203 Segment
X33203 N33203 N33204 Segment
X33204 N33204 N33205 Segment
X33205 N33205 N33206 Segment
X33206 N33206 N33207 Segment
X33207 N33207 N33208 Segment
X33208 N33208 N33209 Segment
X33209 N33209 N33210 Segment
X33210 N33210 N33211 Segment
X33211 N33211 N33212 Segment
X33212 N33212 N33213 Segment
X33213 N33213 N33214 Segment
X33214 N33214 N33215 Segment
X33215 N33215 N33216 Segment
X33216 N33216 N33217 Segment
X33217 N33217 N33218 Segment
X33218 N33218 N33219 Segment
X33219 N33219 N33220 Segment
X33220 N33220 N33221 Segment
X33221 N33221 N33222 Segment
X33222 N33222 N33223 Segment
X33223 N33223 N33224 Segment
X33224 N33224 N33225 Segment
X33225 N33225 N33226 Segment
X33226 N33226 N33227 Segment
X33227 N33227 N33228 Segment
X33228 N33228 N33229 Segment
X33229 N33229 N33230 Segment
X33230 N33230 N33231 Segment
X33231 N33231 N33232 Segment
X33232 N33232 N33233 Segment
X33233 N33233 N33234 Segment
X33234 N33234 N33235 Segment
X33235 N33235 N33236 Segment
X33236 N33236 N33237 Segment
X33237 N33237 N33238 Segment
X33238 N33238 N33239 Segment
X33239 N33239 N33240 Segment
X33240 N33240 N33241 Segment
X33241 N33241 N33242 Segment
X33242 N33242 N33243 Segment
X33243 N33243 N33244 Segment
X33244 N33244 N33245 Segment
X33245 N33245 N33246 Segment
X33246 N33246 N33247 Segment
X33247 N33247 N33248 Segment
X33248 N33248 N33249 Segment
X33249 N33249 N33250 Segment
X33250 N33250 N33251 Segment
X33251 N33251 N33252 Segment
X33252 N33252 N33253 Segment
X33253 N33253 N33254 Segment
X33254 N33254 N33255 Segment
X33255 N33255 N33256 Segment
X33256 N33256 N33257 Segment
X33257 N33257 N33258 Segment
X33258 N33258 N33259 Segment
X33259 N33259 N33260 Segment
X33260 N33260 N33261 Segment
X33261 N33261 N33262 Segment
X33262 N33262 N33263 Segment
X33263 N33263 N33264 Segment
X33264 N33264 N33265 Segment
X33265 N33265 N33266 Segment
X33266 N33266 N33267 Segment
X33267 N33267 N33268 Segment
X33268 N33268 N33269 Segment
X33269 N33269 N33270 Segment
X33270 N33270 N33271 Segment
X33271 N33271 N33272 Segment
X33272 N33272 N33273 Segment
X33273 N33273 N33274 Segment
X33274 N33274 N33275 Segment
X33275 N33275 N33276 Segment
X33276 N33276 N33277 Segment
X33277 N33277 N33278 Segment
X33278 N33278 N33279 Segment
X33279 N33279 N33280 Segment
X33280 N33280 N33281 Segment
X33281 N33281 N33282 Segment
X33282 N33282 N33283 Segment
X33283 N33283 N33284 Segment
X33284 N33284 N33285 Segment
X33285 N33285 N33286 Segment
X33286 N33286 N33287 Segment
X33287 N33287 N33288 Segment
X33288 N33288 N33289 Segment
X33289 N33289 N33290 Segment
X33290 N33290 N33291 Segment
X33291 N33291 N33292 Segment
X33292 N33292 N33293 Segment
X33293 N33293 N33294 Segment
X33294 N33294 N33295 Segment
X33295 N33295 N33296 Segment
X33296 N33296 N33297 Segment
X33297 N33297 N33298 Segment
X33298 N33298 N33299 Segment
X33299 N33299 N33300 Segment
X33300 N33300 N33301 Segment
X33301 N33301 N33302 Segment
X33302 N33302 N33303 Segment
X33303 N33303 N33304 Segment
X33304 N33304 N33305 Segment
X33305 N33305 N33306 Segment
X33306 N33306 N33307 Segment
X33307 N33307 N33308 Segment
X33308 N33308 N33309 Segment
X33309 N33309 N33310 Segment
X33310 N33310 N33311 Segment
X33311 N33311 N33312 Segment
X33312 N33312 N33313 Segment
X33313 N33313 N33314 Segment
X33314 N33314 N33315 Segment
X33315 N33315 N33316 Segment
X33316 N33316 N33317 Segment
X33317 N33317 N33318 Segment
X33318 N33318 N33319 Segment
X33319 N33319 N33320 Segment
X33320 N33320 N33321 Segment
X33321 N33321 N33322 Segment
X33322 N33322 N33323 Segment
X33323 N33323 N33324 Segment
X33324 N33324 N33325 Segment
X33325 N33325 N33326 Segment
X33326 N33326 N33327 Segment
X33327 N33327 N33328 Segment
X33328 N33328 N33329 Segment
X33329 N33329 N33330 Segment
X33330 N33330 N33331 Segment
X33331 N33331 N33332 Segment
X33332 N33332 N33333 Segment
X33333 N33333 N33334 Segment
X33334 N33334 N33335 Segment
X33335 N33335 N33336 Segment
X33336 N33336 N33337 Segment
X33337 N33337 N33338 Segment
X33338 N33338 N33339 Segment
X33339 N33339 N33340 Segment
X33340 N33340 N33341 Segment
X33341 N33341 N33342 Segment
X33342 N33342 N33343 Segment
X33343 N33343 N33344 Segment
X33344 N33344 N33345 Segment
X33345 N33345 N33346 Segment
X33346 N33346 N33347 Segment
X33347 N33347 N33348 Segment
X33348 N33348 N33349 Segment
X33349 N33349 N33350 Segment
X33350 N33350 N33351 Segment
X33351 N33351 N33352 Segment
X33352 N33352 N33353 Segment
X33353 N33353 N33354 Segment
X33354 N33354 N33355 Segment
X33355 N33355 N33356 Segment
X33356 N33356 N33357 Segment
X33357 N33357 N33358 Segment
X33358 N33358 N33359 Segment
X33359 N33359 N33360 Segment
X33360 N33360 N33361 Segment
X33361 N33361 N33362 Segment
X33362 N33362 N33363 Segment
X33363 N33363 N33364 Segment
X33364 N33364 N33365 Segment
X33365 N33365 N33366 Segment
X33366 N33366 N33367 Segment
X33367 N33367 N33368 Segment
X33368 N33368 N33369 Segment
X33369 N33369 N33370 Segment
X33370 N33370 N33371 Segment
X33371 N33371 N33372 Segment
X33372 N33372 N33373 Segment
X33373 N33373 N33374 Segment
X33374 N33374 N33375 Segment
X33375 N33375 N33376 Segment
X33376 N33376 N33377 Segment
X33377 N33377 N33378 Segment
X33378 N33378 N33379 Segment
X33379 N33379 N33380 Segment
X33380 N33380 N33381 Segment
X33381 N33381 N33382 Segment
X33382 N33382 N33383 Segment
X33383 N33383 N33384 Segment
X33384 N33384 N33385 Segment
X33385 N33385 N33386 Segment
X33386 N33386 N33387 Segment
X33387 N33387 N33388 Segment
X33388 N33388 N33389 Segment
X33389 N33389 N33390 Segment
X33390 N33390 N33391 Segment
X33391 N33391 N33392 Segment
X33392 N33392 N33393 Segment
X33393 N33393 N33394 Segment
X33394 N33394 N33395 Segment
X33395 N33395 N33396 Segment
X33396 N33396 N33397 Segment
X33397 N33397 N33398 Segment
X33398 N33398 N33399 Segment
X33399 N33399 N33400 Segment
X33400 N33400 N33401 Segment
X33401 N33401 N33402 Segment
X33402 N33402 N33403 Segment
X33403 N33403 N33404 Segment
X33404 N33404 N33405 Segment
X33405 N33405 N33406 Segment
X33406 N33406 N33407 Segment
X33407 N33407 N33408 Segment
X33408 N33408 N33409 Segment
X33409 N33409 N33410 Segment
X33410 N33410 N33411 Segment
X33411 N33411 N33412 Segment
X33412 N33412 N33413 Segment
X33413 N33413 N33414 Segment
X33414 N33414 N33415 Segment
X33415 N33415 N33416 Segment
X33416 N33416 N33417 Segment
X33417 N33417 N33418 Segment
X33418 N33418 N33419 Segment
X33419 N33419 N33420 Segment
X33420 N33420 N33421 Segment
X33421 N33421 N33422 Segment
X33422 N33422 N33423 Segment
X33423 N33423 N33424 Segment
X33424 N33424 N33425 Segment
X33425 N33425 N33426 Segment
X33426 N33426 N33427 Segment
X33427 N33427 N33428 Segment
X33428 N33428 N33429 Segment
X33429 N33429 N33430 Segment
X33430 N33430 N33431 Segment
X33431 N33431 N33432 Segment
X33432 N33432 N33433 Segment
X33433 N33433 N33434 Segment
X33434 N33434 N33435 Segment
X33435 N33435 N33436 Segment
X33436 N33436 N33437 Segment
X33437 N33437 N33438 Segment
X33438 N33438 N33439 Segment
X33439 N33439 N33440 Segment
X33440 N33440 N33441 Segment
X33441 N33441 N33442 Segment
X33442 N33442 N33443 Segment
X33443 N33443 N33444 Segment
X33444 N33444 N33445 Segment
X33445 N33445 N33446 Segment
X33446 N33446 N33447 Segment
X33447 N33447 N33448 Segment
X33448 N33448 N33449 Segment
X33449 N33449 N33450 Segment
X33450 N33450 N33451 Segment
X33451 N33451 N33452 Segment
X33452 N33452 N33453 Segment
X33453 N33453 N33454 Segment
X33454 N33454 N33455 Segment
X33455 N33455 N33456 Segment
X33456 N33456 N33457 Segment
X33457 N33457 N33458 Segment
X33458 N33458 N33459 Segment
X33459 N33459 N33460 Segment
X33460 N33460 N33461 Segment
X33461 N33461 N33462 Segment
X33462 N33462 N33463 Segment
X33463 N33463 N33464 Segment
X33464 N33464 N33465 Segment
X33465 N33465 N33466 Segment
X33466 N33466 N33467 Segment
X33467 N33467 N33468 Segment
X33468 N33468 N33469 Segment
X33469 N33469 N33470 Segment
X33470 N33470 N33471 Segment
X33471 N33471 N33472 Segment
X33472 N33472 N33473 Segment
X33473 N33473 N33474 Segment
X33474 N33474 N33475 Segment
X33475 N33475 N33476 Segment
X33476 N33476 N33477 Segment
X33477 N33477 N33478 Segment
X33478 N33478 N33479 Segment
X33479 N33479 N33480 Segment
X33480 N33480 N33481 Segment
X33481 N33481 N33482 Segment
X33482 N33482 N33483 Segment
X33483 N33483 N33484 Segment
X33484 N33484 N33485 Segment
X33485 N33485 N33486 Segment
X33486 N33486 N33487 Segment
X33487 N33487 N33488 Segment
X33488 N33488 N33489 Segment
X33489 N33489 N33490 Segment
X33490 N33490 N33491 Segment
X33491 N33491 N33492 Segment
X33492 N33492 N33493 Segment
X33493 N33493 N33494 Segment
X33494 N33494 N33495 Segment
X33495 N33495 N33496 Segment
X33496 N33496 N33497 Segment
X33497 N33497 N33498 Segment
X33498 N33498 N33499 Segment
X33499 N33499 N33500 Segment
X33500 N33500 N33501 Segment
X33501 N33501 N33502 Segment
X33502 N33502 N33503 Segment
X33503 N33503 N33504 Segment
X33504 N33504 N33505 Segment
X33505 N33505 N33506 Segment
X33506 N33506 N33507 Segment
X33507 N33507 N33508 Segment
X33508 N33508 N33509 Segment
X33509 N33509 N33510 Segment
X33510 N33510 N33511 Segment
X33511 N33511 N33512 Segment
X33512 N33512 N33513 Segment
X33513 N33513 N33514 Segment
X33514 N33514 N33515 Segment
X33515 N33515 N33516 Segment
X33516 N33516 N33517 Segment
X33517 N33517 N33518 Segment
X33518 N33518 N33519 Segment
X33519 N33519 N33520 Segment
X33520 N33520 N33521 Segment
X33521 N33521 N33522 Segment
X33522 N33522 N33523 Segment
X33523 N33523 N33524 Segment
X33524 N33524 N33525 Segment
X33525 N33525 N33526 Segment
X33526 N33526 N33527 Segment
X33527 N33527 N33528 Segment
X33528 N33528 N33529 Segment
X33529 N33529 N33530 Segment
X33530 N33530 N33531 Segment
X33531 N33531 N33532 Segment
X33532 N33532 N33533 Segment
X33533 N33533 N33534 Segment
X33534 N33534 N33535 Segment
X33535 N33535 N33536 Segment
X33536 N33536 N33537 Segment
X33537 N33537 N33538 Segment
X33538 N33538 N33539 Segment
X33539 N33539 N33540 Segment
X33540 N33540 N33541 Segment
X33541 N33541 N33542 Segment
X33542 N33542 N33543 Segment
X33543 N33543 N33544 Segment
X33544 N33544 N33545 Segment
X33545 N33545 N33546 Segment
X33546 N33546 N33547 Segment
X33547 N33547 N33548 Segment
X33548 N33548 N33549 Segment
X33549 N33549 N33550 Segment
X33550 N33550 N33551 Segment
X33551 N33551 N33552 Segment
X33552 N33552 N33553 Segment
X33553 N33553 N33554 Segment
X33554 N33554 N33555 Segment
X33555 N33555 N33556 Segment
X33556 N33556 N33557 Segment
X33557 N33557 N33558 Segment
X33558 N33558 N33559 Segment
X33559 N33559 N33560 Segment
X33560 N33560 N33561 Segment
X33561 N33561 N33562 Segment
X33562 N33562 N33563 Segment
X33563 N33563 N33564 Segment
X33564 N33564 N33565 Segment
X33565 N33565 N33566 Segment
X33566 N33566 N33567 Segment
X33567 N33567 N33568 Segment
X33568 N33568 N33569 Segment
X33569 N33569 N33570 Segment
X33570 N33570 N33571 Segment
X33571 N33571 N33572 Segment
X33572 N33572 N33573 Segment
X33573 N33573 N33574 Segment
X33574 N33574 N33575 Segment
X33575 N33575 N33576 Segment
X33576 N33576 N33577 Segment
X33577 N33577 N33578 Segment
X33578 N33578 N33579 Segment
X33579 N33579 N33580 Segment
X33580 N33580 N33581 Segment
X33581 N33581 N33582 Segment
X33582 N33582 N33583 Segment
X33583 N33583 N33584 Segment
X33584 N33584 N33585 Segment
X33585 N33585 N33586 Segment
X33586 N33586 N33587 Segment
X33587 N33587 N33588 Segment
X33588 N33588 N33589 Segment
X33589 N33589 N33590 Segment
X33590 N33590 N33591 Segment
X33591 N33591 N33592 Segment
X33592 N33592 N33593 Segment
X33593 N33593 N33594 Segment
X33594 N33594 N33595 Segment
X33595 N33595 N33596 Segment
X33596 N33596 N33597 Segment
X33597 N33597 N33598 Segment
X33598 N33598 N33599 Segment
X33599 N33599 N33600 Segment
X33600 N33600 N33601 Segment
X33601 N33601 N33602 Segment
X33602 N33602 N33603 Segment
X33603 N33603 N33604 Segment
X33604 N33604 N33605 Segment
X33605 N33605 N33606 Segment
X33606 N33606 N33607 Segment
X33607 N33607 N33608 Segment
X33608 N33608 N33609 Segment
X33609 N33609 N33610 Segment
X33610 N33610 N33611 Segment
X33611 N33611 N33612 Segment
X33612 N33612 N33613 Segment
X33613 N33613 N33614 Segment
X33614 N33614 N33615 Segment
X33615 N33615 N33616 Segment
X33616 N33616 N33617 Segment
X33617 N33617 N33618 Segment
X33618 N33618 N33619 Segment
X33619 N33619 N33620 Segment
X33620 N33620 N33621 Segment
X33621 N33621 N33622 Segment
X33622 N33622 N33623 Segment
X33623 N33623 N33624 Segment
X33624 N33624 N33625 Segment
X33625 N33625 N33626 Segment
X33626 N33626 N33627 Segment
X33627 N33627 N33628 Segment
X33628 N33628 N33629 Segment
X33629 N33629 N33630 Segment
X33630 N33630 N33631 Segment
X33631 N33631 N33632 Segment
X33632 N33632 N33633 Segment
X33633 N33633 N33634 Segment
X33634 N33634 N33635 Segment
X33635 N33635 N33636 Segment
X33636 N33636 N33637 Segment
X33637 N33637 N33638 Segment
X33638 N33638 N33639 Segment
X33639 N33639 N33640 Segment
X33640 N33640 N33641 Segment
X33641 N33641 N33642 Segment
X33642 N33642 N33643 Segment
X33643 N33643 N33644 Segment
X33644 N33644 N33645 Segment
X33645 N33645 N33646 Segment
X33646 N33646 N33647 Segment
X33647 N33647 N33648 Segment
X33648 N33648 N33649 Segment
X33649 N33649 N33650 Segment
X33650 N33650 N33651 Segment
X33651 N33651 N33652 Segment
X33652 N33652 N33653 Segment
X33653 N33653 N33654 Segment
X33654 N33654 N33655 Segment
X33655 N33655 N33656 Segment
X33656 N33656 N33657 Segment
X33657 N33657 N33658 Segment
X33658 N33658 N33659 Segment
X33659 N33659 N33660 Segment
X33660 N33660 N33661 Segment
X33661 N33661 N33662 Segment
X33662 N33662 N33663 Segment
X33663 N33663 N33664 Segment
X33664 N33664 N33665 Segment
X33665 N33665 N33666 Segment
X33666 N33666 N33667 Segment
X33667 N33667 N33668 Segment
X33668 N33668 N33669 Segment
X33669 N33669 N33670 Segment
X33670 N33670 N33671 Segment
X33671 N33671 N33672 Segment
X33672 N33672 N33673 Segment
X33673 N33673 N33674 Segment
X33674 N33674 N33675 Segment
X33675 N33675 N33676 Segment
X33676 N33676 N33677 Segment
X33677 N33677 N33678 Segment
X33678 N33678 N33679 Segment
X33679 N33679 N33680 Segment
X33680 N33680 N33681 Segment
X33681 N33681 N33682 Segment
X33682 N33682 N33683 Segment
X33683 N33683 N33684 Segment
X33684 N33684 N33685 Segment
X33685 N33685 N33686 Segment
X33686 N33686 N33687 Segment
X33687 N33687 N33688 Segment
X33688 N33688 N33689 Segment
X33689 N33689 N33690 Segment
X33690 N33690 N33691 Segment
X33691 N33691 N33692 Segment
X33692 N33692 N33693 Segment
X33693 N33693 N33694 Segment
X33694 N33694 N33695 Segment
X33695 N33695 N33696 Segment
X33696 N33696 N33697 Segment
X33697 N33697 N33698 Segment
X33698 N33698 N33699 Segment
X33699 N33699 N33700 Segment
X33700 N33700 N33701 Segment
X33701 N33701 N33702 Segment
X33702 N33702 N33703 Segment
X33703 N33703 N33704 Segment
X33704 N33704 N33705 Segment
X33705 N33705 N33706 Segment
X33706 N33706 N33707 Segment
X33707 N33707 N33708 Segment
X33708 N33708 N33709 Segment
X33709 N33709 N33710 Segment
X33710 N33710 N33711 Segment
X33711 N33711 N33712 Segment
X33712 N33712 N33713 Segment
X33713 N33713 N33714 Segment
X33714 N33714 N33715 Segment
X33715 N33715 N33716 Segment
X33716 N33716 N33717 Segment
X33717 N33717 N33718 Segment
X33718 N33718 N33719 Segment
X33719 N33719 N33720 Segment
X33720 N33720 N33721 Segment
X33721 N33721 N33722 Segment
X33722 N33722 N33723 Segment
X33723 N33723 N33724 Segment
X33724 N33724 N33725 Segment
X33725 N33725 N33726 Segment
X33726 N33726 N33727 Segment
X33727 N33727 N33728 Segment
X33728 N33728 N33729 Segment
X33729 N33729 N33730 Segment
X33730 N33730 N33731 Segment
X33731 N33731 N33732 Segment
X33732 N33732 N33733 Segment
X33733 N33733 N33734 Segment
X33734 N33734 N33735 Segment
X33735 N33735 N33736 Segment
X33736 N33736 N33737 Segment
X33737 N33737 N33738 Segment
X33738 N33738 N33739 Segment
X33739 N33739 N33740 Segment
X33740 N33740 N33741 Segment
X33741 N33741 N33742 Segment
X33742 N33742 N33743 Segment
X33743 N33743 N33744 Segment
X33744 N33744 N33745 Segment
X33745 N33745 N33746 Segment
X33746 N33746 N33747 Segment
X33747 N33747 N33748 Segment
X33748 N33748 N33749 Segment
X33749 N33749 N33750 Segment
X33750 N33750 N33751 Segment
X33751 N33751 N33752 Segment
X33752 N33752 N33753 Segment
X33753 N33753 N33754 Segment
X33754 N33754 N33755 Segment
X33755 N33755 N33756 Segment
X33756 N33756 N33757 Segment
X33757 N33757 N33758 Segment
X33758 N33758 N33759 Segment
X33759 N33759 N33760 Segment
X33760 N33760 N33761 Segment
X33761 N33761 N33762 Segment
X33762 N33762 N33763 Segment
X33763 N33763 N33764 Segment
X33764 N33764 N33765 Segment
X33765 N33765 N33766 Segment
X33766 N33766 N33767 Segment
X33767 N33767 N33768 Segment
X33768 N33768 N33769 Segment
X33769 N33769 N33770 Segment
X33770 N33770 N33771 Segment
X33771 N33771 N33772 Segment
X33772 N33772 N33773 Segment
X33773 N33773 N33774 Segment
X33774 N33774 N33775 Segment
X33775 N33775 N33776 Segment
X33776 N33776 N33777 Segment
X33777 N33777 N33778 Segment
X33778 N33778 N33779 Segment
X33779 N33779 N33780 Segment
X33780 N33780 N33781 Segment
X33781 N33781 N33782 Segment
X33782 N33782 N33783 Segment
X33783 N33783 N33784 Segment
X33784 N33784 N33785 Segment
X33785 N33785 N33786 Segment
X33786 N33786 N33787 Segment
X33787 N33787 N33788 Segment
X33788 N33788 N33789 Segment
X33789 N33789 N33790 Segment
X33790 N33790 N33791 Segment
X33791 N33791 N33792 Segment
X33792 N33792 N33793 Segment
X33793 N33793 N33794 Segment
X33794 N33794 N33795 Segment
X33795 N33795 N33796 Segment
X33796 N33796 N33797 Segment
X33797 N33797 N33798 Segment
X33798 N33798 N33799 Segment
X33799 N33799 N33800 Segment
X33800 N33800 N33801 Segment
X33801 N33801 N33802 Segment
X33802 N33802 N33803 Segment
X33803 N33803 N33804 Segment
X33804 N33804 N33805 Segment
X33805 N33805 N33806 Segment
X33806 N33806 N33807 Segment
X33807 N33807 N33808 Segment
X33808 N33808 N33809 Segment
X33809 N33809 N33810 Segment
X33810 N33810 N33811 Segment
X33811 N33811 N33812 Segment
X33812 N33812 N33813 Segment
X33813 N33813 N33814 Segment
X33814 N33814 N33815 Segment
X33815 N33815 N33816 Segment
X33816 N33816 N33817 Segment
X33817 N33817 N33818 Segment
X33818 N33818 N33819 Segment
X33819 N33819 N33820 Segment
X33820 N33820 N33821 Segment
X33821 N33821 N33822 Segment
X33822 N33822 N33823 Segment
X33823 N33823 N33824 Segment
X33824 N33824 N33825 Segment
X33825 N33825 N33826 Segment
X33826 N33826 N33827 Segment
X33827 N33827 N33828 Segment
X33828 N33828 N33829 Segment
X33829 N33829 N33830 Segment
X33830 N33830 N33831 Segment
X33831 N33831 N33832 Segment
X33832 N33832 N33833 Segment
X33833 N33833 N33834 Segment
X33834 N33834 N33835 Segment
X33835 N33835 N33836 Segment
X33836 N33836 N33837 Segment
X33837 N33837 N33838 Segment
X33838 N33838 N33839 Segment
X33839 N33839 N33840 Segment
X33840 N33840 N33841 Segment
X33841 N33841 N33842 Segment
X33842 N33842 N33843 Segment
X33843 N33843 N33844 Segment
X33844 N33844 N33845 Segment
X33845 N33845 N33846 Segment
X33846 N33846 N33847 Segment
X33847 N33847 N33848 Segment
X33848 N33848 N33849 Segment
X33849 N33849 N33850 Segment
X33850 N33850 N33851 Segment
X33851 N33851 N33852 Segment
X33852 N33852 N33853 Segment
X33853 N33853 N33854 Segment
X33854 N33854 N33855 Segment
X33855 N33855 N33856 Segment
X33856 N33856 N33857 Segment
X33857 N33857 N33858 Segment
X33858 N33858 N33859 Segment
X33859 N33859 N33860 Segment
X33860 N33860 N33861 Segment
X33861 N33861 N33862 Segment
X33862 N33862 N33863 Segment
X33863 N33863 N33864 Segment
X33864 N33864 N33865 Segment
X33865 N33865 N33866 Segment
X33866 N33866 N33867 Segment
X33867 N33867 N33868 Segment
X33868 N33868 N33869 Segment
X33869 N33869 N33870 Segment
X33870 N33870 N33871 Segment
X33871 N33871 N33872 Segment
X33872 N33872 N33873 Segment
X33873 N33873 N33874 Segment
X33874 N33874 N33875 Segment
X33875 N33875 N33876 Segment
X33876 N33876 N33877 Segment
X33877 N33877 N33878 Segment
X33878 N33878 N33879 Segment
X33879 N33879 N33880 Segment
X33880 N33880 N33881 Segment
X33881 N33881 N33882 Segment
X33882 N33882 N33883 Segment
X33883 N33883 N33884 Segment
X33884 N33884 N33885 Segment
X33885 N33885 N33886 Segment
X33886 N33886 N33887 Segment
X33887 N33887 N33888 Segment
X33888 N33888 N33889 Segment
X33889 N33889 N33890 Segment
X33890 N33890 N33891 Segment
X33891 N33891 N33892 Segment
X33892 N33892 N33893 Segment
X33893 N33893 N33894 Segment
X33894 N33894 N33895 Segment
X33895 N33895 N33896 Segment
X33896 N33896 N33897 Segment
X33897 N33897 N33898 Segment
X33898 N33898 N33899 Segment
X33899 N33899 N33900 Segment
X33900 N33900 N33901 Segment
X33901 N33901 N33902 Segment
X33902 N33902 N33903 Segment
X33903 N33903 N33904 Segment
X33904 N33904 N33905 Segment
X33905 N33905 N33906 Segment
X33906 N33906 N33907 Segment
X33907 N33907 N33908 Segment
X33908 N33908 N33909 Segment
X33909 N33909 N33910 Segment
X33910 N33910 N33911 Segment
X33911 N33911 N33912 Segment
X33912 N33912 N33913 Segment
X33913 N33913 N33914 Segment
X33914 N33914 N33915 Segment
X33915 N33915 N33916 Segment
X33916 N33916 N33917 Segment
X33917 N33917 N33918 Segment
X33918 N33918 N33919 Segment
X33919 N33919 N33920 Segment
X33920 N33920 N33921 Segment
X33921 N33921 N33922 Segment
X33922 N33922 N33923 Segment
X33923 N33923 N33924 Segment
X33924 N33924 N33925 Segment
X33925 N33925 N33926 Segment
X33926 N33926 N33927 Segment
X33927 N33927 N33928 Segment
X33928 N33928 N33929 Segment
X33929 N33929 N33930 Segment
X33930 N33930 N33931 Segment
X33931 N33931 N33932 Segment
X33932 N33932 N33933 Segment
X33933 N33933 N33934 Segment
X33934 N33934 N33935 Segment
X33935 N33935 N33936 Segment
X33936 N33936 N33937 Segment
X33937 N33937 N33938 Segment
X33938 N33938 N33939 Segment
X33939 N33939 N33940 Segment
X33940 N33940 N33941 Segment
X33941 N33941 N33942 Segment
X33942 N33942 N33943 Segment
X33943 N33943 N33944 Segment
X33944 N33944 N33945 Segment
X33945 N33945 N33946 Segment
X33946 N33946 N33947 Segment
X33947 N33947 N33948 Segment
X33948 N33948 N33949 Segment
X33949 N33949 N33950 Segment
X33950 N33950 N33951 Segment
X33951 N33951 N33952 Segment
X33952 N33952 N33953 Segment
X33953 N33953 N33954 Segment
X33954 N33954 N33955 Segment
X33955 N33955 N33956 Segment
X33956 N33956 N33957 Segment
X33957 N33957 N33958 Segment
X33958 N33958 N33959 Segment
X33959 N33959 N33960 Segment
X33960 N33960 N33961 Segment
X33961 N33961 N33962 Segment
X33962 N33962 N33963 Segment
X33963 N33963 N33964 Segment
X33964 N33964 N33965 Segment
X33965 N33965 N33966 Segment
X33966 N33966 N33967 Segment
X33967 N33967 N33968 Segment
X33968 N33968 N33969 Segment
X33969 N33969 N33970 Segment
X33970 N33970 N33971 Segment
X33971 N33971 N33972 Segment
X33972 N33972 N33973 Segment
X33973 N33973 N33974 Segment
X33974 N33974 N33975 Segment
X33975 N33975 N33976 Segment
X33976 N33976 N33977 Segment
X33977 N33977 N33978 Segment
X33978 N33978 N33979 Segment
X33979 N33979 N33980 Segment
X33980 N33980 N33981 Segment
X33981 N33981 N33982 Segment
X33982 N33982 N33983 Segment
X33983 N33983 N33984 Segment
X33984 N33984 N33985 Segment
X33985 N33985 N33986 Segment
X33986 N33986 N33987 Segment
X33987 N33987 N33988 Segment
X33988 N33988 N33989 Segment
X33989 N33989 N33990 Segment
X33990 N33990 N33991 Segment
X33991 N33991 N33992 Segment
X33992 N33992 N33993 Segment
X33993 N33993 N33994 Segment
X33994 N33994 N33995 Segment
X33995 N33995 N33996 Segment
X33996 N33996 N33997 Segment
X33997 N33997 N33998 Segment
X33998 N33998 N33999 Segment
X33999 N33999 N34000 Segment
X34000 N34000 N34001 Segment
X34001 N34001 N34002 Segment
X34002 N34002 N34003 Segment
X34003 N34003 N34004 Segment
X34004 N34004 N34005 Segment
X34005 N34005 N34006 Segment
X34006 N34006 N34007 Segment
X34007 N34007 N34008 Segment
X34008 N34008 N34009 Segment
X34009 N34009 N34010 Segment
X34010 N34010 N34011 Segment
X34011 N34011 N34012 Segment
X34012 N34012 N34013 Segment
X34013 N34013 N34014 Segment
X34014 N34014 N34015 Segment
X34015 N34015 N34016 Segment
X34016 N34016 N34017 Segment
X34017 N34017 N34018 Segment
X34018 N34018 N34019 Segment
X34019 N34019 N34020 Segment
X34020 N34020 N34021 Segment
X34021 N34021 N34022 Segment
X34022 N34022 N34023 Segment
X34023 N34023 N34024 Segment
X34024 N34024 N34025 Segment
X34025 N34025 N34026 Segment
X34026 N34026 N34027 Segment
X34027 N34027 N34028 Segment
X34028 N34028 N34029 Segment
X34029 N34029 N34030 Segment
X34030 N34030 N34031 Segment
X34031 N34031 N34032 Segment
X34032 N34032 N34033 Segment
X34033 N34033 N34034 Segment
X34034 N34034 N34035 Segment
X34035 N34035 N34036 Segment
X34036 N34036 N34037 Segment
X34037 N34037 N34038 Segment
X34038 N34038 N34039 Segment
X34039 N34039 N34040 Segment
X34040 N34040 N34041 Segment
X34041 N34041 N34042 Segment
X34042 N34042 N34043 Segment
X34043 N34043 N34044 Segment
X34044 N34044 N34045 Segment
X34045 N34045 N34046 Segment
X34046 N34046 N34047 Segment
X34047 N34047 N34048 Segment
X34048 N34048 N34049 Segment
X34049 N34049 N34050 Segment
X34050 N34050 N34051 Segment
X34051 N34051 N34052 Segment
X34052 N34052 N34053 Segment
X34053 N34053 N34054 Segment
X34054 N34054 N34055 Segment
X34055 N34055 N34056 Segment
X34056 N34056 N34057 Segment
X34057 N34057 N34058 Segment
X34058 N34058 N34059 Segment
X34059 N34059 N34060 Segment
X34060 N34060 N34061 Segment
X34061 N34061 N34062 Segment
X34062 N34062 N34063 Segment
X34063 N34063 N34064 Segment
X34064 N34064 N34065 Segment
X34065 N34065 N34066 Segment
X34066 N34066 N34067 Segment
X34067 N34067 N34068 Segment
X34068 N34068 N34069 Segment
X34069 N34069 N34070 Segment
X34070 N34070 N34071 Segment
X34071 N34071 N34072 Segment
X34072 N34072 N34073 Segment
X34073 N34073 N34074 Segment
X34074 N34074 N34075 Segment
X34075 N34075 N34076 Segment
X34076 N34076 N34077 Segment
X34077 N34077 N34078 Segment
X34078 N34078 N34079 Segment
X34079 N34079 N34080 Segment
X34080 N34080 N34081 Segment
X34081 N34081 N34082 Segment
X34082 N34082 N34083 Segment
X34083 N34083 N34084 Segment
X34084 N34084 N34085 Segment
X34085 N34085 N34086 Segment
X34086 N34086 N34087 Segment
X34087 N34087 N34088 Segment
X34088 N34088 N34089 Segment
X34089 N34089 N34090 Segment
X34090 N34090 N34091 Segment
X34091 N34091 N34092 Segment
X34092 N34092 N34093 Segment
X34093 N34093 N34094 Segment
X34094 N34094 N34095 Segment
X34095 N34095 N34096 Segment
X34096 N34096 N34097 Segment
X34097 N34097 N34098 Segment
X34098 N34098 N34099 Segment
X34099 N34099 N34100 Segment
X34100 N34100 N34101 Segment
X34101 N34101 N34102 Segment
X34102 N34102 N34103 Segment
X34103 N34103 N34104 Segment
X34104 N34104 N34105 Segment
X34105 N34105 N34106 Segment
X34106 N34106 N34107 Segment
X34107 N34107 N34108 Segment
X34108 N34108 N34109 Segment
X34109 N34109 N34110 Segment
X34110 N34110 N34111 Segment
X34111 N34111 N34112 Segment
X34112 N34112 N34113 Segment
X34113 N34113 N34114 Segment
X34114 N34114 N34115 Segment
X34115 N34115 N34116 Segment
X34116 N34116 N34117 Segment
X34117 N34117 N34118 Segment
X34118 N34118 N34119 Segment
X34119 N34119 N34120 Segment
X34120 N34120 N34121 Segment
X34121 N34121 N34122 Segment
X34122 N34122 N34123 Segment
X34123 N34123 N34124 Segment
X34124 N34124 N34125 Segment
X34125 N34125 N34126 Segment
X34126 N34126 N34127 Segment
X34127 N34127 N34128 Segment
X34128 N34128 N34129 Segment
X34129 N34129 N34130 Segment
X34130 N34130 N34131 Segment
X34131 N34131 N34132 Segment
X34132 N34132 N34133 Segment
X34133 N34133 N34134 Segment
X34134 N34134 N34135 Segment
X34135 N34135 N34136 Segment
X34136 N34136 N34137 Segment
X34137 N34137 N34138 Segment
X34138 N34138 N34139 Segment
X34139 N34139 N34140 Segment
X34140 N34140 N34141 Segment
X34141 N34141 N34142 Segment
X34142 N34142 N34143 Segment
X34143 N34143 N34144 Segment
X34144 N34144 N34145 Segment
X34145 N34145 N34146 Segment
X34146 N34146 N34147 Segment
X34147 N34147 N34148 Segment
X34148 N34148 N34149 Segment
X34149 N34149 N34150 Segment
X34150 N34150 N34151 Segment
X34151 N34151 N34152 Segment
X34152 N34152 N34153 Segment
X34153 N34153 N34154 Segment
X34154 N34154 N34155 Segment
X34155 N34155 N34156 Segment
X34156 N34156 N34157 Segment
X34157 N34157 N34158 Segment
X34158 N34158 N34159 Segment
X34159 N34159 N34160 Segment
X34160 N34160 N34161 Segment
X34161 N34161 N34162 Segment
X34162 N34162 N34163 Segment
X34163 N34163 N34164 Segment
X34164 N34164 N34165 Segment
X34165 N34165 N34166 Segment
X34166 N34166 N34167 Segment
X34167 N34167 N34168 Segment
X34168 N34168 N34169 Segment
X34169 N34169 N34170 Segment
X34170 N34170 N34171 Segment
X34171 N34171 N34172 Segment
X34172 N34172 N34173 Segment
X34173 N34173 N34174 Segment
X34174 N34174 N34175 Segment
X34175 N34175 N34176 Segment
X34176 N34176 N34177 Segment
X34177 N34177 N34178 Segment
X34178 N34178 N34179 Segment
X34179 N34179 N34180 Segment
X34180 N34180 N34181 Segment
X34181 N34181 N34182 Segment
X34182 N34182 N34183 Segment
X34183 N34183 N34184 Segment
X34184 N34184 N34185 Segment
X34185 N34185 N34186 Segment
X34186 N34186 N34187 Segment
X34187 N34187 N34188 Segment
X34188 N34188 N34189 Segment
X34189 N34189 N34190 Segment
X34190 N34190 N34191 Segment
X34191 N34191 N34192 Segment
X34192 N34192 N34193 Segment
X34193 N34193 N34194 Segment
X34194 N34194 N34195 Segment
X34195 N34195 N34196 Segment
X34196 N34196 N34197 Segment
X34197 N34197 N34198 Segment
X34198 N34198 N34199 Segment
X34199 N34199 N34200 Segment
X34200 N34200 N34201 Segment
X34201 N34201 N34202 Segment
X34202 N34202 N34203 Segment
X34203 N34203 N34204 Segment
X34204 N34204 N34205 Segment
X34205 N34205 N34206 Segment
X34206 N34206 N34207 Segment
X34207 N34207 N34208 Segment
X34208 N34208 N34209 Segment
X34209 N34209 N34210 Segment
X34210 N34210 N34211 Segment
X34211 N34211 N34212 Segment
X34212 N34212 N34213 Segment
X34213 N34213 N34214 Segment
X34214 N34214 N34215 Segment
X34215 N34215 N34216 Segment
X34216 N34216 N34217 Segment
X34217 N34217 N34218 Segment
X34218 N34218 N34219 Segment
X34219 N34219 N34220 Segment
X34220 N34220 N34221 Segment
X34221 N34221 N34222 Segment
X34222 N34222 N34223 Segment
X34223 N34223 N34224 Segment
X34224 N34224 N34225 Segment
X34225 N34225 N34226 Segment
X34226 N34226 N34227 Segment
X34227 N34227 N34228 Segment
X34228 N34228 N34229 Segment
X34229 N34229 N34230 Segment
X34230 N34230 N34231 Segment
X34231 N34231 N34232 Segment
X34232 N34232 N34233 Segment
X34233 N34233 N34234 Segment
X34234 N34234 N34235 Segment
X34235 N34235 N34236 Segment
X34236 N34236 N34237 Segment
X34237 N34237 N34238 Segment
X34238 N34238 N34239 Segment
X34239 N34239 N34240 Segment
X34240 N34240 N34241 Segment
X34241 N34241 N34242 Segment
X34242 N34242 N34243 Segment
X34243 N34243 N34244 Segment
X34244 N34244 N34245 Segment
X34245 N34245 N34246 Segment
X34246 N34246 N34247 Segment
X34247 N34247 N34248 Segment
X34248 N34248 N34249 Segment
X34249 N34249 N34250 Segment
X34250 N34250 N34251 Segment
X34251 N34251 N34252 Segment
X34252 N34252 N34253 Segment
X34253 N34253 N34254 Segment
X34254 N34254 N34255 Segment
X34255 N34255 N34256 Segment
X34256 N34256 N34257 Segment
X34257 N34257 N34258 Segment
X34258 N34258 N34259 Segment
X34259 N34259 N34260 Segment
X34260 N34260 N34261 Segment
X34261 N34261 N34262 Segment
X34262 N34262 N34263 Segment
X34263 N34263 N34264 Segment
X34264 N34264 N34265 Segment
X34265 N34265 N34266 Segment
X34266 N34266 N34267 Segment
X34267 N34267 N34268 Segment
X34268 N34268 N34269 Segment
X34269 N34269 N34270 Segment
X34270 N34270 N34271 Segment
X34271 N34271 N34272 Segment
X34272 N34272 N34273 Segment
X34273 N34273 N34274 Segment
X34274 N34274 N34275 Segment
X34275 N34275 N34276 Segment
X34276 N34276 N34277 Segment
X34277 N34277 N34278 Segment
X34278 N34278 N34279 Segment
X34279 N34279 N34280 Segment
X34280 N34280 N34281 Segment
X34281 N34281 N34282 Segment
X34282 N34282 N34283 Segment
X34283 N34283 N34284 Segment
X34284 N34284 N34285 Segment
X34285 N34285 N34286 Segment
X34286 N34286 N34287 Segment
X34287 N34287 N34288 Segment
X34288 N34288 N34289 Segment
X34289 N34289 N34290 Segment
X34290 N34290 N34291 Segment
X34291 N34291 N34292 Segment
X34292 N34292 N34293 Segment
X34293 N34293 N34294 Segment
X34294 N34294 N34295 Segment
X34295 N34295 N34296 Segment
X34296 N34296 N34297 Segment
X34297 N34297 N34298 Segment
X34298 N34298 N34299 Segment
X34299 N34299 N34300 Segment
X34300 N34300 N34301 Segment
X34301 N34301 N34302 Segment
X34302 N34302 N34303 Segment
X34303 N34303 N34304 Segment
X34304 N34304 N34305 Segment
X34305 N34305 N34306 Segment
X34306 N34306 N34307 Segment
X34307 N34307 N34308 Segment
X34308 N34308 N34309 Segment
X34309 N34309 N34310 Segment
X34310 N34310 N34311 Segment
X34311 N34311 N34312 Segment
X34312 N34312 N34313 Segment
X34313 N34313 N34314 Segment
X34314 N34314 N34315 Segment
X34315 N34315 N34316 Segment
X34316 N34316 N34317 Segment
X34317 N34317 N34318 Segment
X34318 N34318 N34319 Segment
X34319 N34319 N34320 Segment
X34320 N34320 N34321 Segment
X34321 N34321 N34322 Segment
X34322 N34322 N34323 Segment
X34323 N34323 N34324 Segment
X34324 N34324 N34325 Segment
X34325 N34325 N34326 Segment
X34326 N34326 N34327 Segment
X34327 N34327 N34328 Segment
X34328 N34328 N34329 Segment
X34329 N34329 N34330 Segment
X34330 N34330 N34331 Segment
X34331 N34331 N34332 Segment
X34332 N34332 N34333 Segment
X34333 N34333 N34334 Segment
X34334 N34334 N34335 Segment
X34335 N34335 N34336 Segment
X34336 N34336 N34337 Segment
X34337 N34337 N34338 Segment
X34338 N34338 N34339 Segment
X34339 N34339 N34340 Segment
X34340 N34340 N34341 Segment
X34341 N34341 N34342 Segment
X34342 N34342 N34343 Segment
X34343 N34343 N34344 Segment
X34344 N34344 N34345 Segment
X34345 N34345 N34346 Segment
X34346 N34346 N34347 Segment
X34347 N34347 N34348 Segment
X34348 N34348 N34349 Segment
X34349 N34349 N34350 Segment
X34350 N34350 N34351 Segment
X34351 N34351 N34352 Segment
X34352 N34352 N34353 Segment
X34353 N34353 N34354 Segment
X34354 N34354 N34355 Segment
X34355 N34355 N34356 Segment
X34356 N34356 N34357 Segment
X34357 N34357 N34358 Segment
X34358 N34358 N34359 Segment
X34359 N34359 N34360 Segment
X34360 N34360 N34361 Segment
X34361 N34361 N34362 Segment
X34362 N34362 N34363 Segment
X34363 N34363 N34364 Segment
X34364 N34364 N34365 Segment
X34365 N34365 N34366 Segment
X34366 N34366 N34367 Segment
X34367 N34367 N34368 Segment
X34368 N34368 N34369 Segment
X34369 N34369 N34370 Segment
X34370 N34370 N34371 Segment
X34371 N34371 N34372 Segment
X34372 N34372 N34373 Segment
X34373 N34373 N34374 Segment
X34374 N34374 N34375 Segment
X34375 N34375 N34376 Segment
X34376 N34376 N34377 Segment
X34377 N34377 N34378 Segment
X34378 N34378 N34379 Segment
X34379 N34379 N34380 Segment
X34380 N34380 N34381 Segment
X34381 N34381 N34382 Segment
X34382 N34382 N34383 Segment
X34383 N34383 N34384 Segment
X34384 N34384 N34385 Segment
X34385 N34385 N34386 Segment
X34386 N34386 N34387 Segment
X34387 N34387 N34388 Segment
X34388 N34388 N34389 Segment
X34389 N34389 N34390 Segment
X34390 N34390 N34391 Segment
X34391 N34391 N34392 Segment
X34392 N34392 N34393 Segment
X34393 N34393 N34394 Segment
X34394 N34394 N34395 Segment
X34395 N34395 N34396 Segment
X34396 N34396 N34397 Segment
X34397 N34397 N34398 Segment
X34398 N34398 N34399 Segment
X34399 N34399 N34400 Segment
X34400 N34400 N34401 Segment
X34401 N34401 N34402 Segment
X34402 N34402 N34403 Segment
X34403 N34403 N34404 Segment
X34404 N34404 N34405 Segment
X34405 N34405 N34406 Segment
X34406 N34406 N34407 Segment
X34407 N34407 N34408 Segment
X34408 N34408 N34409 Segment
X34409 N34409 N34410 Segment
X34410 N34410 N34411 Segment
X34411 N34411 N34412 Segment
X34412 N34412 N34413 Segment
X34413 N34413 N34414 Segment
X34414 N34414 N34415 Segment
X34415 N34415 N34416 Segment
X34416 N34416 N34417 Segment
X34417 N34417 N34418 Segment
X34418 N34418 N34419 Segment
X34419 N34419 N34420 Segment
X34420 N34420 N34421 Segment
X34421 N34421 N34422 Segment
X34422 N34422 N34423 Segment
X34423 N34423 N34424 Segment
X34424 N34424 N34425 Segment
X34425 N34425 N34426 Segment
X34426 N34426 N34427 Segment
X34427 N34427 N34428 Segment
X34428 N34428 N34429 Segment
X34429 N34429 N34430 Segment
X34430 N34430 N34431 Segment
X34431 N34431 N34432 Segment
X34432 N34432 N34433 Segment
X34433 N34433 N34434 Segment
X34434 N34434 N34435 Segment
X34435 N34435 N34436 Segment
X34436 N34436 N34437 Segment
X34437 N34437 N34438 Segment
X34438 N34438 N34439 Segment
X34439 N34439 N34440 Segment
X34440 N34440 N34441 Segment
X34441 N34441 N34442 Segment
X34442 N34442 N34443 Segment
X34443 N34443 N34444 Segment
X34444 N34444 N34445 Segment
X34445 N34445 N34446 Segment
X34446 N34446 N34447 Segment
X34447 N34447 N34448 Segment
X34448 N34448 N34449 Segment
X34449 N34449 N34450 Segment
X34450 N34450 N34451 Segment
X34451 N34451 N34452 Segment
X34452 N34452 N34453 Segment
X34453 N34453 N34454 Segment
X34454 N34454 N34455 Segment
X34455 N34455 N34456 Segment
X34456 N34456 N34457 Segment
X34457 N34457 N34458 Segment
X34458 N34458 N34459 Segment
X34459 N34459 N34460 Segment
X34460 N34460 N34461 Segment
X34461 N34461 N34462 Segment
X34462 N34462 N34463 Segment
X34463 N34463 N34464 Segment
X34464 N34464 N34465 Segment
X34465 N34465 N34466 Segment
X34466 N34466 N34467 Segment
X34467 N34467 N34468 Segment
X34468 N34468 N34469 Segment
X34469 N34469 N34470 Segment
X34470 N34470 N34471 Segment
X34471 N34471 N34472 Segment
X34472 N34472 N34473 Segment
X34473 N34473 N34474 Segment
X34474 N34474 N34475 Segment
X34475 N34475 N34476 Segment
X34476 N34476 N34477 Segment
X34477 N34477 N34478 Segment
X34478 N34478 N34479 Segment
X34479 N34479 N34480 Segment
X34480 N34480 N34481 Segment
X34481 N34481 N34482 Segment
X34482 N34482 N34483 Segment
X34483 N34483 N34484 Segment
X34484 N34484 N34485 Segment
X34485 N34485 N34486 Segment
X34486 N34486 N34487 Segment
X34487 N34487 N34488 Segment
X34488 N34488 N34489 Segment
X34489 N34489 N34490 Segment
X34490 N34490 N34491 Segment
X34491 N34491 N34492 Segment
X34492 N34492 N34493 Segment
X34493 N34493 N34494 Segment
X34494 N34494 N34495 Segment
X34495 N34495 N34496 Segment
X34496 N34496 N34497 Segment
X34497 N34497 N34498 Segment
X34498 N34498 N34499 Segment
X34499 N34499 N34500 Segment
X34500 N34500 N34501 Segment
X34501 N34501 N34502 Segment
X34502 N34502 N34503 Segment
X34503 N34503 N34504 Segment
X34504 N34504 N34505 Segment
X34505 N34505 N34506 Segment
X34506 N34506 N34507 Segment
X34507 N34507 N34508 Segment
X34508 N34508 N34509 Segment
X34509 N34509 N34510 Segment
X34510 N34510 N34511 Segment
X34511 N34511 N34512 Segment
X34512 N34512 N34513 Segment
X34513 N34513 N34514 Segment
X34514 N34514 N34515 Segment
X34515 N34515 N34516 Segment
X34516 N34516 N34517 Segment
X34517 N34517 N34518 Segment
X34518 N34518 N34519 Segment
X34519 N34519 N34520 Segment
X34520 N34520 N34521 Segment
X34521 N34521 N34522 Segment
X34522 N34522 N34523 Segment
X34523 N34523 N34524 Segment
X34524 N34524 N34525 Segment
X34525 N34525 N34526 Segment
X34526 N34526 N34527 Segment
X34527 N34527 N34528 Segment
X34528 N34528 N34529 Segment
X34529 N34529 N34530 Segment
X34530 N34530 N34531 Segment
X34531 N34531 N34532 Segment
X34532 N34532 N34533 Segment
X34533 N34533 N34534 Segment
X34534 N34534 N34535 Segment
X34535 N34535 N34536 Segment
X34536 N34536 N34537 Segment
X34537 N34537 N34538 Segment
X34538 N34538 N34539 Segment
X34539 N34539 N34540 Segment
X34540 N34540 N34541 Segment
X34541 N34541 N34542 Segment
X34542 N34542 N34543 Segment
X34543 N34543 N34544 Segment
X34544 N34544 N34545 Segment
X34545 N34545 N34546 Segment
X34546 N34546 N34547 Segment
X34547 N34547 N34548 Segment
X34548 N34548 N34549 Segment
X34549 N34549 N34550 Segment
X34550 N34550 N34551 Segment
X34551 N34551 N34552 Segment
X34552 N34552 N34553 Segment
X34553 N34553 N34554 Segment
X34554 N34554 N34555 Segment
X34555 N34555 N34556 Segment
X34556 N34556 N34557 Segment
X34557 N34557 N34558 Segment
X34558 N34558 N34559 Segment
X34559 N34559 N34560 Segment
X34560 N34560 N34561 Segment
X34561 N34561 N34562 Segment
X34562 N34562 N34563 Segment
X34563 N34563 N34564 Segment
X34564 N34564 N34565 Segment
X34565 N34565 N34566 Segment
X34566 N34566 N34567 Segment
X34567 N34567 N34568 Segment
X34568 N34568 N34569 Segment
X34569 N34569 N34570 Segment
X34570 N34570 N34571 Segment
X34571 N34571 N34572 Segment
X34572 N34572 N34573 Segment
X34573 N34573 N34574 Segment
X34574 N34574 N34575 Segment
X34575 N34575 N34576 Segment
X34576 N34576 N34577 Segment
X34577 N34577 N34578 Segment
X34578 N34578 N34579 Segment
X34579 N34579 N34580 Segment
X34580 N34580 N34581 Segment
X34581 N34581 N34582 Segment
X34582 N34582 N34583 Segment
X34583 N34583 N34584 Segment
X34584 N34584 N34585 Segment
X34585 N34585 N34586 Segment
X34586 N34586 N34587 Segment
X34587 N34587 N34588 Segment
X34588 N34588 N34589 Segment
X34589 N34589 N34590 Segment
X34590 N34590 N34591 Segment
X34591 N34591 N34592 Segment
X34592 N34592 N34593 Segment
X34593 N34593 N34594 Segment
X34594 N34594 N34595 Segment
X34595 N34595 N34596 Segment
X34596 N34596 N34597 Segment
X34597 N34597 N34598 Segment
X34598 N34598 N34599 Segment
X34599 N34599 N34600 Segment
X34600 N34600 N34601 Segment
X34601 N34601 N34602 Segment
X34602 N34602 N34603 Segment
X34603 N34603 N34604 Segment
X34604 N34604 N34605 Segment
X34605 N34605 N34606 Segment
X34606 N34606 N34607 Segment
X34607 N34607 N34608 Segment
X34608 N34608 N34609 Segment
X34609 N34609 N34610 Segment
X34610 N34610 N34611 Segment
X34611 N34611 N34612 Segment
X34612 N34612 N34613 Segment
X34613 N34613 N34614 Segment
X34614 N34614 N34615 Segment
X34615 N34615 N34616 Segment
X34616 N34616 N34617 Segment
X34617 N34617 N34618 Segment
X34618 N34618 N34619 Segment
X34619 N34619 N34620 Segment
X34620 N34620 N34621 Segment
X34621 N34621 N34622 Segment
X34622 N34622 N34623 Segment
X34623 N34623 N34624 Segment
X34624 N34624 N34625 Segment
X34625 N34625 N34626 Segment
X34626 N34626 N34627 Segment
X34627 N34627 N34628 Segment
X34628 N34628 N34629 Segment
X34629 N34629 N34630 Segment
X34630 N34630 N34631 Segment
X34631 N34631 N34632 Segment
X34632 N34632 N34633 Segment
X34633 N34633 N34634 Segment
X34634 N34634 N34635 Segment
X34635 N34635 N34636 Segment
X34636 N34636 N34637 Segment
X34637 N34637 N34638 Segment
X34638 N34638 N34639 Segment
X34639 N34639 N34640 Segment
X34640 N34640 N34641 Segment
X34641 N34641 N34642 Segment
X34642 N34642 N34643 Segment
X34643 N34643 N34644 Segment
X34644 N34644 N34645 Segment
X34645 N34645 N34646 Segment
X34646 N34646 N34647 Segment
X34647 N34647 N34648 Segment
X34648 N34648 N34649 Segment
X34649 N34649 N34650 Segment
X34650 N34650 N34651 Segment
X34651 N34651 N34652 Segment
X34652 N34652 N34653 Segment
X34653 N34653 N34654 Segment
X34654 N34654 N34655 Segment
X34655 N34655 N34656 Segment
X34656 N34656 N34657 Segment
X34657 N34657 N34658 Segment
X34658 N34658 N34659 Segment
X34659 N34659 N34660 Segment
X34660 N34660 N34661 Segment
X34661 N34661 N34662 Segment
X34662 N34662 N34663 Segment
X34663 N34663 N34664 Segment
X34664 N34664 N34665 Segment
X34665 N34665 N34666 Segment
X34666 N34666 N34667 Segment
X34667 N34667 N34668 Segment
X34668 N34668 N34669 Segment
X34669 N34669 N34670 Segment
X34670 N34670 N34671 Segment
X34671 N34671 N34672 Segment
X34672 N34672 N34673 Segment
X34673 N34673 N34674 Segment
X34674 N34674 N34675 Segment
X34675 N34675 N34676 Segment
X34676 N34676 N34677 Segment
X34677 N34677 N34678 Segment
X34678 N34678 N34679 Segment
X34679 N34679 N34680 Segment
X34680 N34680 N34681 Segment
X34681 N34681 N34682 Segment
X34682 N34682 N34683 Segment
X34683 N34683 N34684 Segment
X34684 N34684 N34685 Segment
X34685 N34685 N34686 Segment
X34686 N34686 N34687 Segment
X34687 N34687 N34688 Segment
X34688 N34688 N34689 Segment
X34689 N34689 N34690 Segment
X34690 N34690 N34691 Segment
X34691 N34691 N34692 Segment
X34692 N34692 N34693 Segment
X34693 N34693 N34694 Segment
X34694 N34694 N34695 Segment
X34695 N34695 N34696 Segment
X34696 N34696 N34697 Segment
X34697 N34697 N34698 Segment
X34698 N34698 N34699 Segment
X34699 N34699 N34700 Segment
X34700 N34700 N34701 Segment
X34701 N34701 N34702 Segment
X34702 N34702 N34703 Segment
X34703 N34703 N34704 Segment
X34704 N34704 N34705 Segment
X34705 N34705 N34706 Segment
X34706 N34706 N34707 Segment
X34707 N34707 N34708 Segment
X34708 N34708 N34709 Segment
X34709 N34709 N34710 Segment
X34710 N34710 N34711 Segment
X34711 N34711 N34712 Segment
X34712 N34712 N34713 Segment
X34713 N34713 N34714 Segment
X34714 N34714 N34715 Segment
X34715 N34715 N34716 Segment
X34716 N34716 N34717 Segment
X34717 N34717 N34718 Segment
X34718 N34718 N34719 Segment
X34719 N34719 N34720 Segment
X34720 N34720 N34721 Segment
X34721 N34721 N34722 Segment
X34722 N34722 N34723 Segment
X34723 N34723 N34724 Segment
X34724 N34724 N34725 Segment
X34725 N34725 N34726 Segment
X34726 N34726 N34727 Segment
X34727 N34727 N34728 Segment
X34728 N34728 N34729 Segment
X34729 N34729 N34730 Segment
X34730 N34730 N34731 Segment
X34731 N34731 N34732 Segment
X34732 N34732 N34733 Segment
X34733 N34733 N34734 Segment
X34734 N34734 N34735 Segment
X34735 N34735 N34736 Segment
X34736 N34736 N34737 Segment
X34737 N34737 N34738 Segment
X34738 N34738 N34739 Segment
X34739 N34739 N34740 Segment
X34740 N34740 N34741 Segment
X34741 N34741 N34742 Segment
X34742 N34742 N34743 Segment
X34743 N34743 N34744 Segment
X34744 N34744 N34745 Segment
X34745 N34745 N34746 Segment
X34746 N34746 N34747 Segment
X34747 N34747 N34748 Segment
X34748 N34748 N34749 Segment
X34749 N34749 N34750 Segment
X34750 N34750 N34751 Segment
X34751 N34751 N34752 Segment
X34752 N34752 N34753 Segment
X34753 N34753 N34754 Segment
X34754 N34754 N34755 Segment
X34755 N34755 N34756 Segment
X34756 N34756 N34757 Segment
X34757 N34757 N34758 Segment
X34758 N34758 N34759 Segment
X34759 N34759 N34760 Segment
X34760 N34760 N34761 Segment
X34761 N34761 N34762 Segment
X34762 N34762 N34763 Segment
X34763 N34763 N34764 Segment
X34764 N34764 N34765 Segment
X34765 N34765 N34766 Segment
X34766 N34766 N34767 Segment
X34767 N34767 N34768 Segment
X34768 N34768 N34769 Segment
X34769 N34769 N34770 Segment
X34770 N34770 N34771 Segment
X34771 N34771 N34772 Segment
X34772 N34772 N34773 Segment
X34773 N34773 N34774 Segment
X34774 N34774 N34775 Segment
X34775 N34775 N34776 Segment
X34776 N34776 N34777 Segment
X34777 N34777 N34778 Segment
X34778 N34778 N34779 Segment
X34779 N34779 N34780 Segment
X34780 N34780 N34781 Segment
X34781 N34781 N34782 Segment
X34782 N34782 N34783 Segment
X34783 N34783 N34784 Segment
X34784 N34784 N34785 Segment
X34785 N34785 N34786 Segment
X34786 N34786 N34787 Segment
X34787 N34787 N34788 Segment
X34788 N34788 N34789 Segment
X34789 N34789 N34790 Segment
X34790 N34790 N34791 Segment
X34791 N34791 N34792 Segment
X34792 N34792 N34793 Segment
X34793 N34793 N34794 Segment
X34794 N34794 N34795 Segment
X34795 N34795 N34796 Segment
X34796 N34796 N34797 Segment
X34797 N34797 N34798 Segment
X34798 N34798 N34799 Segment
X34799 N34799 N34800 Segment
X34800 N34800 N34801 Segment
X34801 N34801 N34802 Segment
X34802 N34802 N34803 Segment
X34803 N34803 N34804 Segment
X34804 N34804 N34805 Segment
X34805 N34805 N34806 Segment
X34806 N34806 N34807 Segment
X34807 N34807 N34808 Segment
X34808 N34808 N34809 Segment
X34809 N34809 N34810 Segment
X34810 N34810 N34811 Segment
X34811 N34811 N34812 Segment
X34812 N34812 N34813 Segment
X34813 N34813 N34814 Segment
X34814 N34814 N34815 Segment
X34815 N34815 N34816 Segment
X34816 N34816 N34817 Segment
X34817 N34817 N34818 Segment
X34818 N34818 N34819 Segment
X34819 N34819 N34820 Segment
X34820 N34820 N34821 Segment
X34821 N34821 N34822 Segment
X34822 N34822 N34823 Segment
X34823 N34823 N34824 Segment
X34824 N34824 N34825 Segment
X34825 N34825 N34826 Segment
X34826 N34826 N34827 Segment
X34827 N34827 N34828 Segment
X34828 N34828 N34829 Segment
X34829 N34829 N34830 Segment
X34830 N34830 N34831 Segment
X34831 N34831 N34832 Segment
X34832 N34832 N34833 Segment
X34833 N34833 N34834 Segment
X34834 N34834 N34835 Segment
X34835 N34835 N34836 Segment
X34836 N34836 N34837 Segment
X34837 N34837 N34838 Segment
X34838 N34838 N34839 Segment
X34839 N34839 N34840 Segment
X34840 N34840 N34841 Segment
X34841 N34841 N34842 Segment
X34842 N34842 N34843 Segment
X34843 N34843 N34844 Segment
X34844 N34844 N34845 Segment
X34845 N34845 N34846 Segment
X34846 N34846 N34847 Segment
X34847 N34847 N34848 Segment
X34848 N34848 N34849 Segment
X34849 N34849 N34850 Segment
X34850 N34850 N34851 Segment
X34851 N34851 N34852 Segment
X34852 N34852 N34853 Segment
X34853 N34853 N34854 Segment
X34854 N34854 N34855 Segment
X34855 N34855 N34856 Segment
X34856 N34856 N34857 Segment
X34857 N34857 N34858 Segment
X34858 N34858 N34859 Segment
X34859 N34859 N34860 Segment
X34860 N34860 N34861 Segment
X34861 N34861 N34862 Segment
X34862 N34862 N34863 Segment
X34863 N34863 N34864 Segment
X34864 N34864 N34865 Segment
X34865 N34865 N34866 Segment
X34866 N34866 N34867 Segment
X34867 N34867 N34868 Segment
X34868 N34868 N34869 Segment
X34869 N34869 N34870 Segment
X34870 N34870 N34871 Segment
X34871 N34871 N34872 Segment
X34872 N34872 N34873 Segment
X34873 N34873 N34874 Segment
X34874 N34874 N34875 Segment
X34875 N34875 N34876 Segment
X34876 N34876 N34877 Segment
X34877 N34877 N34878 Segment
X34878 N34878 N34879 Segment
X34879 N34879 N34880 Segment
X34880 N34880 N34881 Segment
X34881 N34881 N34882 Segment
X34882 N34882 N34883 Segment
X34883 N34883 N34884 Segment
X34884 N34884 N34885 Segment
X34885 N34885 N34886 Segment
X34886 N34886 N34887 Segment
X34887 N34887 N34888 Segment
X34888 N34888 N34889 Segment
X34889 N34889 N34890 Segment
X34890 N34890 N34891 Segment
X34891 N34891 N34892 Segment
X34892 N34892 N34893 Segment
X34893 N34893 N34894 Segment
X34894 N34894 N34895 Segment
X34895 N34895 N34896 Segment
X34896 N34896 N34897 Segment
X34897 N34897 N34898 Segment
X34898 N34898 N34899 Segment
X34899 N34899 N34900 Segment
X34900 N34900 N34901 Segment
X34901 N34901 N34902 Segment
X34902 N34902 N34903 Segment
X34903 N34903 N34904 Segment
X34904 N34904 N34905 Segment
X34905 N34905 N34906 Segment
X34906 N34906 N34907 Segment
X34907 N34907 N34908 Segment
X34908 N34908 N34909 Segment
X34909 N34909 N34910 Segment
X34910 N34910 N34911 Segment
X34911 N34911 N34912 Segment
X34912 N34912 N34913 Segment
X34913 N34913 N34914 Segment
X34914 N34914 N34915 Segment
X34915 N34915 N34916 Segment
X34916 N34916 N34917 Segment
X34917 N34917 N34918 Segment
X34918 N34918 N34919 Segment
X34919 N34919 N34920 Segment
X34920 N34920 N34921 Segment
X34921 N34921 N34922 Segment
X34922 N34922 N34923 Segment
X34923 N34923 N34924 Segment
X34924 N34924 N34925 Segment
X34925 N34925 N34926 Segment
X34926 N34926 N34927 Segment
X34927 N34927 N34928 Segment
X34928 N34928 N34929 Segment
X34929 N34929 N34930 Segment
X34930 N34930 N34931 Segment
X34931 N34931 N34932 Segment
X34932 N34932 N34933 Segment
X34933 N34933 N34934 Segment
X34934 N34934 N34935 Segment
X34935 N34935 N34936 Segment
X34936 N34936 N34937 Segment
X34937 N34937 N34938 Segment
X34938 N34938 N34939 Segment
X34939 N34939 N34940 Segment
X34940 N34940 N34941 Segment
X34941 N34941 N34942 Segment
X34942 N34942 N34943 Segment
X34943 N34943 N34944 Segment
X34944 N34944 N34945 Segment
X34945 N34945 N34946 Segment
X34946 N34946 N34947 Segment
X34947 N34947 N34948 Segment
X34948 N34948 N34949 Segment
X34949 N34949 N34950 Segment
X34950 N34950 N34951 Segment
X34951 N34951 N34952 Segment
X34952 N34952 N34953 Segment
X34953 N34953 N34954 Segment
X34954 N34954 N34955 Segment
X34955 N34955 N34956 Segment
X34956 N34956 N34957 Segment
X34957 N34957 N34958 Segment
X34958 N34958 N34959 Segment
X34959 N34959 N34960 Segment
X34960 N34960 N34961 Segment
X34961 N34961 N34962 Segment
X34962 N34962 N34963 Segment
X34963 N34963 N34964 Segment
X34964 N34964 N34965 Segment
X34965 N34965 N34966 Segment
X34966 N34966 N34967 Segment
X34967 N34967 N34968 Segment
X34968 N34968 N34969 Segment
X34969 N34969 N34970 Segment
X34970 N34970 N34971 Segment
X34971 N34971 N34972 Segment
X34972 N34972 N34973 Segment
X34973 N34973 N34974 Segment
X34974 N34974 N34975 Segment
X34975 N34975 N34976 Segment
X34976 N34976 N34977 Segment
X34977 N34977 N34978 Segment
X34978 N34978 N34979 Segment
X34979 N34979 N34980 Segment
X34980 N34980 N34981 Segment
X34981 N34981 N34982 Segment
X34982 N34982 N34983 Segment
X34983 N34983 N34984 Segment
X34984 N34984 N34985 Segment
X34985 N34985 N34986 Segment
X34986 N34986 N34987 Segment
X34987 N34987 N34988 Segment
X34988 N34988 N34989 Segment
X34989 N34989 N34990 Segment
X34990 N34990 N34991 Segment
X34991 N34991 N34992 Segment
X34992 N34992 N34993 Segment
X34993 N34993 N34994 Segment
X34994 N34994 N34995 Segment
X34995 N34995 N34996 Segment
X34996 N34996 N34997 Segment
X34997 N34997 N34998 Segment
X34998 N34998 N34999 Segment
X34999 N34999 N35000 Segment
X35000 N35000 N35001 Segment
X35001 N35001 N35002 Segment
X35002 N35002 N35003 Segment
X35003 N35003 N35004 Segment
X35004 N35004 N35005 Segment
X35005 N35005 N35006 Segment
X35006 N35006 N35007 Segment
X35007 N35007 N35008 Segment
X35008 N35008 N35009 Segment
X35009 N35009 N35010 Segment
X35010 N35010 N35011 Segment
X35011 N35011 N35012 Segment
X35012 N35012 N35013 Segment
X35013 N35013 N35014 Segment
X35014 N35014 N35015 Segment
X35015 N35015 N35016 Segment
X35016 N35016 N35017 Segment
X35017 N35017 N35018 Segment
X35018 N35018 N35019 Segment
X35019 N35019 N35020 Segment
X35020 N35020 N35021 Segment
X35021 N35021 N35022 Segment
X35022 N35022 N35023 Segment
X35023 N35023 N35024 Segment
X35024 N35024 N35025 Segment
X35025 N35025 N35026 Segment
X35026 N35026 N35027 Segment
X35027 N35027 N35028 Segment
X35028 N35028 N35029 Segment
X35029 N35029 N35030 Segment
X35030 N35030 N35031 Segment
X35031 N35031 N35032 Segment
X35032 N35032 N35033 Segment
X35033 N35033 N35034 Segment
X35034 N35034 N35035 Segment
X35035 N35035 N35036 Segment
X35036 N35036 N35037 Segment
X35037 N35037 N35038 Segment
X35038 N35038 N35039 Segment
X35039 N35039 N35040 Segment
X35040 N35040 N35041 Segment
X35041 N35041 N35042 Segment
X35042 N35042 N35043 Segment
X35043 N35043 N35044 Segment
X35044 N35044 N35045 Segment
X35045 N35045 N35046 Segment
X35046 N35046 N35047 Segment
X35047 N35047 N35048 Segment
X35048 N35048 N35049 Segment
X35049 N35049 N35050 Segment
X35050 N35050 N35051 Segment
X35051 N35051 N35052 Segment
X35052 N35052 N35053 Segment
X35053 N35053 N35054 Segment
X35054 N35054 N35055 Segment
X35055 N35055 N35056 Segment
X35056 N35056 N35057 Segment
X35057 N35057 N35058 Segment
X35058 N35058 N35059 Segment
X35059 N35059 N35060 Segment
X35060 N35060 N35061 Segment
X35061 N35061 N35062 Segment
X35062 N35062 N35063 Segment
X35063 N35063 N35064 Segment
X35064 N35064 N35065 Segment
X35065 N35065 N35066 Segment
X35066 N35066 N35067 Segment
X35067 N35067 N35068 Segment
X35068 N35068 N35069 Segment
X35069 N35069 N35070 Segment
X35070 N35070 N35071 Segment
X35071 N35071 N35072 Segment
X35072 N35072 N35073 Segment
X35073 N35073 N35074 Segment
X35074 N35074 N35075 Segment
X35075 N35075 N35076 Segment
X35076 N35076 N35077 Segment
X35077 N35077 N35078 Segment
X35078 N35078 N35079 Segment
X35079 N35079 N35080 Segment
X35080 N35080 N35081 Segment
X35081 N35081 N35082 Segment
X35082 N35082 N35083 Segment
X35083 N35083 N35084 Segment
X35084 N35084 N35085 Segment
X35085 N35085 N35086 Segment
X35086 N35086 N35087 Segment
X35087 N35087 N35088 Segment
X35088 N35088 N35089 Segment
X35089 N35089 N35090 Segment
X35090 N35090 N35091 Segment
X35091 N35091 N35092 Segment
X35092 N35092 N35093 Segment
X35093 N35093 N35094 Segment
X35094 N35094 N35095 Segment
X35095 N35095 N35096 Segment
X35096 N35096 N35097 Segment
X35097 N35097 N35098 Segment
X35098 N35098 N35099 Segment
X35099 N35099 N35100 Segment
X35100 N35100 N35101 Segment
X35101 N35101 N35102 Segment
X35102 N35102 N35103 Segment
X35103 N35103 N35104 Segment
X35104 N35104 N35105 Segment
X35105 N35105 N35106 Segment
X35106 N35106 N35107 Segment
X35107 N35107 N35108 Segment
X35108 N35108 N35109 Segment
X35109 N35109 N35110 Segment
X35110 N35110 N35111 Segment
X35111 N35111 N35112 Segment
X35112 N35112 N35113 Segment
X35113 N35113 N35114 Segment
X35114 N35114 N35115 Segment
X35115 N35115 N35116 Segment
X35116 N35116 N35117 Segment
X35117 N35117 N35118 Segment
X35118 N35118 N35119 Segment
X35119 N35119 N35120 Segment
X35120 N35120 N35121 Segment
X35121 N35121 N35122 Segment
X35122 N35122 N35123 Segment
X35123 N35123 N35124 Segment
X35124 N35124 N35125 Segment
X35125 N35125 N35126 Segment
X35126 N35126 N35127 Segment
X35127 N35127 N35128 Segment
X35128 N35128 N35129 Segment
X35129 N35129 N35130 Segment
X35130 N35130 N35131 Segment
X35131 N35131 N35132 Segment
X35132 N35132 N35133 Segment
X35133 N35133 N35134 Segment
X35134 N35134 N35135 Segment
X35135 N35135 N35136 Segment
X35136 N35136 N35137 Segment
X35137 N35137 N35138 Segment
X35138 N35138 N35139 Segment
X35139 N35139 N35140 Segment
X35140 N35140 N35141 Segment
X35141 N35141 N35142 Segment
X35142 N35142 N35143 Segment
X35143 N35143 N35144 Segment
X35144 N35144 N35145 Segment
X35145 N35145 N35146 Segment
X35146 N35146 N35147 Segment
X35147 N35147 N35148 Segment
X35148 N35148 N35149 Segment
X35149 N35149 N35150 Segment
X35150 N35150 N35151 Segment
X35151 N35151 N35152 Segment
X35152 N35152 N35153 Segment
X35153 N35153 N35154 Segment
X35154 N35154 N35155 Segment
X35155 N35155 N35156 Segment
X35156 N35156 N35157 Segment
X35157 N35157 N35158 Segment
X35158 N35158 N35159 Segment
X35159 N35159 N35160 Segment
X35160 N35160 N35161 Segment
X35161 N35161 N35162 Segment
X35162 N35162 N35163 Segment
X35163 N35163 N35164 Segment
X35164 N35164 N35165 Segment
X35165 N35165 N35166 Segment
X35166 N35166 N35167 Segment
X35167 N35167 N35168 Segment
X35168 N35168 N35169 Segment
X35169 N35169 N35170 Segment
X35170 N35170 N35171 Segment
X35171 N35171 N35172 Segment
X35172 N35172 N35173 Segment
X35173 N35173 N35174 Segment
X35174 N35174 N35175 Segment
X35175 N35175 N35176 Segment
X35176 N35176 N35177 Segment
X35177 N35177 N35178 Segment
X35178 N35178 N35179 Segment
X35179 N35179 N35180 Segment
X35180 N35180 N35181 Segment
X35181 N35181 N35182 Segment
X35182 N35182 N35183 Segment
X35183 N35183 N35184 Segment
X35184 N35184 N35185 Segment
X35185 N35185 N35186 Segment
X35186 N35186 N35187 Segment
X35187 N35187 N35188 Segment
X35188 N35188 N35189 Segment
X35189 N35189 N35190 Segment
X35190 N35190 N35191 Segment
X35191 N35191 N35192 Segment
X35192 N35192 N35193 Segment
X35193 N35193 N35194 Segment
X35194 N35194 N35195 Segment
X35195 N35195 N35196 Segment
X35196 N35196 N35197 Segment
X35197 N35197 N35198 Segment
X35198 N35198 N35199 Segment
X35199 N35199 N35200 Segment
X35200 N35200 N35201 Segment
X35201 N35201 N35202 Segment
X35202 N35202 N35203 Segment
X35203 N35203 N35204 Segment
X35204 N35204 N35205 Segment
X35205 N35205 N35206 Segment
X35206 N35206 N35207 Segment
X35207 N35207 N35208 Segment
X35208 N35208 N35209 Segment
X35209 N35209 N35210 Segment
X35210 N35210 N35211 Segment
X35211 N35211 N35212 Segment
X35212 N35212 N35213 Segment
X35213 N35213 N35214 Segment
X35214 N35214 N35215 Segment
X35215 N35215 N35216 Segment
X35216 N35216 N35217 Segment
X35217 N35217 N35218 Segment
X35218 N35218 N35219 Segment
X35219 N35219 N35220 Segment
X35220 N35220 N35221 Segment
X35221 N35221 N35222 Segment
X35222 N35222 N35223 Segment
X35223 N35223 N35224 Segment
X35224 N35224 N35225 Segment
X35225 N35225 N35226 Segment
X35226 N35226 N35227 Segment
X35227 N35227 N35228 Segment
X35228 N35228 N35229 Segment
X35229 N35229 N35230 Segment
X35230 N35230 N35231 Segment
X35231 N35231 N35232 Segment
X35232 N35232 N35233 Segment
X35233 N35233 N35234 Segment
X35234 N35234 N35235 Segment
X35235 N35235 N35236 Segment
X35236 N35236 N35237 Segment
X35237 N35237 N35238 Segment
X35238 N35238 N35239 Segment
X35239 N35239 N35240 Segment
X35240 N35240 N35241 Segment
X35241 N35241 N35242 Segment
X35242 N35242 N35243 Segment
X35243 N35243 N35244 Segment
X35244 N35244 N35245 Segment
X35245 N35245 N35246 Segment
X35246 N35246 N35247 Segment
X35247 N35247 N35248 Segment
X35248 N35248 N35249 Segment
X35249 N35249 N35250 Segment
X35250 N35250 N35251 Segment
X35251 N35251 N35252 Segment
X35252 N35252 N35253 Segment
X35253 N35253 N35254 Segment
X35254 N35254 N35255 Segment
X35255 N35255 N35256 Segment
X35256 N35256 N35257 Segment
X35257 N35257 N35258 Segment
X35258 N35258 N35259 Segment
X35259 N35259 N35260 Segment
X35260 N35260 N35261 Segment
X35261 N35261 N35262 Segment
X35262 N35262 N35263 Segment
X35263 N35263 N35264 Segment
X35264 N35264 N35265 Segment
X35265 N35265 N35266 Segment
X35266 N35266 N35267 Segment
X35267 N35267 N35268 Segment
X35268 N35268 N35269 Segment
X35269 N35269 N35270 Segment
X35270 N35270 N35271 Segment
X35271 N35271 N35272 Segment
X35272 N35272 N35273 Segment
X35273 N35273 N35274 Segment
X35274 N35274 N35275 Segment
X35275 N35275 N35276 Segment
X35276 N35276 N35277 Segment
X35277 N35277 N35278 Segment
X35278 N35278 N35279 Segment
X35279 N35279 N35280 Segment
X35280 N35280 N35281 Segment
X35281 N35281 N35282 Segment
X35282 N35282 N35283 Segment
X35283 N35283 N35284 Segment
X35284 N35284 N35285 Segment
X35285 N35285 N35286 Segment
X35286 N35286 N35287 Segment
X35287 N35287 N35288 Segment
X35288 N35288 N35289 Segment
X35289 N35289 N35290 Segment
X35290 N35290 N35291 Segment
X35291 N35291 N35292 Segment
X35292 N35292 N35293 Segment
X35293 N35293 N35294 Segment
X35294 N35294 N35295 Segment
X35295 N35295 N35296 Segment
X35296 N35296 N35297 Segment
X35297 N35297 N35298 Segment
X35298 N35298 N35299 Segment
X35299 N35299 N35300 Segment
X35300 N35300 N35301 Segment
X35301 N35301 N35302 Segment
X35302 N35302 N35303 Segment
X35303 N35303 N35304 Segment
X35304 N35304 N35305 Segment
X35305 N35305 N35306 Segment
X35306 N35306 N35307 Segment
X35307 N35307 N35308 Segment
X35308 N35308 N35309 Segment
X35309 N35309 N35310 Segment
X35310 N35310 N35311 Segment
X35311 N35311 N35312 Segment
X35312 N35312 N35313 Segment
X35313 N35313 N35314 Segment
X35314 N35314 N35315 Segment
X35315 N35315 N35316 Segment
X35316 N35316 N35317 Segment
X35317 N35317 N35318 Segment
X35318 N35318 N35319 Segment
X35319 N35319 N35320 Segment
X35320 N35320 N35321 Segment
X35321 N35321 N35322 Segment
X35322 N35322 N35323 Segment
X35323 N35323 N35324 Segment
X35324 N35324 N35325 Segment
X35325 N35325 N35326 Segment
X35326 N35326 N35327 Segment
X35327 N35327 N35328 Segment
X35328 N35328 N35329 Segment
X35329 N35329 N35330 Segment
X35330 N35330 N35331 Segment
X35331 N35331 N35332 Segment
X35332 N35332 N35333 Segment
X35333 N35333 N35334 Segment
X35334 N35334 N35335 Segment
X35335 N35335 N35336 Segment
X35336 N35336 N35337 Segment
X35337 N35337 N35338 Segment
X35338 N35338 N35339 Segment
X35339 N35339 N35340 Segment
X35340 N35340 N35341 Segment
X35341 N35341 N35342 Segment
X35342 N35342 N35343 Segment
X35343 N35343 N35344 Segment
X35344 N35344 N35345 Segment
X35345 N35345 N35346 Segment
X35346 N35346 N35347 Segment
X35347 N35347 N35348 Segment
X35348 N35348 N35349 Segment
X35349 N35349 N35350 Segment
X35350 N35350 N35351 Segment
X35351 N35351 N35352 Segment
X35352 N35352 N35353 Segment
X35353 N35353 N35354 Segment
X35354 N35354 N35355 Segment
X35355 N35355 N35356 Segment
X35356 N35356 N35357 Segment
X35357 N35357 N35358 Segment
X35358 N35358 N35359 Segment
X35359 N35359 N35360 Segment
X35360 N35360 N35361 Segment
X35361 N35361 N35362 Segment
X35362 N35362 N35363 Segment
X35363 N35363 N35364 Segment
X35364 N35364 N35365 Segment
X35365 N35365 N35366 Segment
X35366 N35366 N35367 Segment
X35367 N35367 N35368 Segment
X35368 N35368 N35369 Segment
X35369 N35369 N35370 Segment
X35370 N35370 N35371 Segment
X35371 N35371 N35372 Segment
X35372 N35372 N35373 Segment
X35373 N35373 N35374 Segment
X35374 N35374 N35375 Segment
X35375 N35375 N35376 Segment
X35376 N35376 N35377 Segment
X35377 N35377 N35378 Segment
X35378 N35378 N35379 Segment
X35379 N35379 N35380 Segment
X35380 N35380 N35381 Segment
X35381 N35381 N35382 Segment
X35382 N35382 N35383 Segment
X35383 N35383 N35384 Segment
X35384 N35384 N35385 Segment
X35385 N35385 N35386 Segment
X35386 N35386 N35387 Segment
X35387 N35387 N35388 Segment
X35388 N35388 N35389 Segment
X35389 N35389 N35390 Segment
X35390 N35390 N35391 Segment
X35391 N35391 N35392 Segment
X35392 N35392 N35393 Segment
X35393 N35393 N35394 Segment
X35394 N35394 N35395 Segment
X35395 N35395 N35396 Segment
X35396 N35396 N35397 Segment
X35397 N35397 N35398 Segment
X35398 N35398 N35399 Segment
X35399 N35399 N35400 Segment
X35400 N35400 N35401 Segment
X35401 N35401 N35402 Segment
X35402 N35402 N35403 Segment
X35403 N35403 N35404 Segment
X35404 N35404 N35405 Segment
X35405 N35405 N35406 Segment
X35406 N35406 N35407 Segment
X35407 N35407 N35408 Segment
X35408 N35408 N35409 Segment
X35409 N35409 N35410 Segment
X35410 N35410 N35411 Segment
X35411 N35411 N35412 Segment
X35412 N35412 N35413 Segment
X35413 N35413 N35414 Segment
X35414 N35414 N35415 Segment
X35415 N35415 N35416 Segment
X35416 N35416 N35417 Segment
X35417 N35417 N35418 Segment
X35418 N35418 N35419 Segment
X35419 N35419 N35420 Segment
X35420 N35420 N35421 Segment
X35421 N35421 N35422 Segment
X35422 N35422 N35423 Segment
X35423 N35423 N35424 Segment
X35424 N35424 N35425 Segment
X35425 N35425 N35426 Segment
X35426 N35426 N35427 Segment
X35427 N35427 N35428 Segment
X35428 N35428 N35429 Segment
X35429 N35429 N35430 Segment
X35430 N35430 N35431 Segment
X35431 N35431 N35432 Segment
X35432 N35432 N35433 Segment
X35433 N35433 N35434 Segment
X35434 N35434 N35435 Segment
X35435 N35435 N35436 Segment
X35436 N35436 N35437 Segment
X35437 N35437 N35438 Segment
X35438 N35438 N35439 Segment
X35439 N35439 N35440 Segment
X35440 N35440 N35441 Segment
X35441 N35441 N35442 Segment
X35442 N35442 N35443 Segment
X35443 N35443 N35444 Segment
X35444 N35444 N35445 Segment
X35445 N35445 N35446 Segment
X35446 N35446 N35447 Segment
X35447 N35447 N35448 Segment
X35448 N35448 N35449 Segment
X35449 N35449 N35450 Segment
X35450 N35450 N35451 Segment
X35451 N35451 N35452 Segment
X35452 N35452 N35453 Segment
X35453 N35453 N35454 Segment
X35454 N35454 N35455 Segment
X35455 N35455 N35456 Segment
X35456 N35456 N35457 Segment
X35457 N35457 N35458 Segment
X35458 N35458 N35459 Segment
X35459 N35459 N35460 Segment
X35460 N35460 N35461 Segment
X35461 N35461 N35462 Segment
X35462 N35462 N35463 Segment
X35463 N35463 N35464 Segment
X35464 N35464 N35465 Segment
X35465 N35465 N35466 Segment
X35466 N35466 N35467 Segment
X35467 N35467 N35468 Segment
X35468 N35468 N35469 Segment
X35469 N35469 N35470 Segment
X35470 N35470 N35471 Segment
X35471 N35471 N35472 Segment
X35472 N35472 N35473 Segment
X35473 N35473 N35474 Segment
X35474 N35474 N35475 Segment
X35475 N35475 N35476 Segment
X35476 N35476 N35477 Segment
X35477 N35477 N35478 Segment
X35478 N35478 N35479 Segment
X35479 N35479 N35480 Segment
X35480 N35480 N35481 Segment
X35481 N35481 N35482 Segment
X35482 N35482 N35483 Segment
X35483 N35483 N35484 Segment
X35484 N35484 N35485 Segment
X35485 N35485 N35486 Segment
X35486 N35486 N35487 Segment
X35487 N35487 N35488 Segment
X35488 N35488 N35489 Segment
X35489 N35489 N35490 Segment
X35490 N35490 N35491 Segment
X35491 N35491 N35492 Segment
X35492 N35492 N35493 Segment
X35493 N35493 N35494 Segment
X35494 N35494 N35495 Segment
X35495 N35495 N35496 Segment
X35496 N35496 N35497 Segment
X35497 N35497 N35498 Segment
X35498 N35498 N35499 Segment
X35499 N35499 N35500 Segment
X35500 N35500 N35501 Segment
X35501 N35501 N35502 Segment
X35502 N35502 N35503 Segment
X35503 N35503 N35504 Segment
X35504 N35504 N35505 Segment
X35505 N35505 N35506 Segment
X35506 N35506 N35507 Segment
X35507 N35507 N35508 Segment
X35508 N35508 N35509 Segment
X35509 N35509 N35510 Segment
X35510 N35510 N35511 Segment
X35511 N35511 N35512 Segment
X35512 N35512 N35513 Segment
X35513 N35513 N35514 Segment
X35514 N35514 N35515 Segment
X35515 N35515 N35516 Segment
X35516 N35516 N35517 Segment
X35517 N35517 N35518 Segment
X35518 N35518 N35519 Segment
X35519 N35519 N35520 Segment
X35520 N35520 N35521 Segment
X35521 N35521 N35522 Segment
X35522 N35522 N35523 Segment
X35523 N35523 N35524 Segment
X35524 N35524 N35525 Segment
X35525 N35525 N35526 Segment
X35526 N35526 N35527 Segment
X35527 N35527 N35528 Segment
X35528 N35528 N35529 Segment
X35529 N35529 N35530 Segment
X35530 N35530 N35531 Segment
X35531 N35531 N35532 Segment
X35532 N35532 N35533 Segment
X35533 N35533 N35534 Segment
X35534 N35534 N35535 Segment
X35535 N35535 N35536 Segment
X35536 N35536 N35537 Segment
X35537 N35537 N35538 Segment
X35538 N35538 N35539 Segment
X35539 N35539 N35540 Segment
X35540 N35540 N35541 Segment
X35541 N35541 N35542 Segment
X35542 N35542 N35543 Segment
X35543 N35543 N35544 Segment
X35544 N35544 N35545 Segment
X35545 N35545 N35546 Segment
X35546 N35546 N35547 Segment
X35547 N35547 N35548 Segment
X35548 N35548 N35549 Segment
X35549 N35549 N35550 Segment
X35550 N35550 N35551 Segment
X35551 N35551 N35552 Segment
X35552 N35552 N35553 Segment
X35553 N35553 N35554 Segment
X35554 N35554 N35555 Segment
X35555 N35555 N35556 Segment
X35556 N35556 N35557 Segment
X35557 N35557 N35558 Segment
X35558 N35558 N35559 Segment
X35559 N35559 N35560 Segment
X35560 N35560 N35561 Segment
X35561 N35561 N35562 Segment
X35562 N35562 N35563 Segment
X35563 N35563 N35564 Segment
X35564 N35564 N35565 Segment
X35565 N35565 N35566 Segment
X35566 N35566 N35567 Segment
X35567 N35567 N35568 Segment
X35568 N35568 N35569 Segment
X35569 N35569 N35570 Segment
X35570 N35570 N35571 Segment
X35571 N35571 N35572 Segment
X35572 N35572 N35573 Segment
X35573 N35573 N35574 Segment
X35574 N35574 N35575 Segment
X35575 N35575 N35576 Segment
X35576 N35576 N35577 Segment
X35577 N35577 N35578 Segment
X35578 N35578 N35579 Segment
X35579 N35579 N35580 Segment
X35580 N35580 N35581 Segment
X35581 N35581 N35582 Segment
X35582 N35582 N35583 Segment
X35583 N35583 N35584 Segment
X35584 N35584 N35585 Segment
X35585 N35585 N35586 Segment
X35586 N35586 N35587 Segment
X35587 N35587 N35588 Segment
X35588 N35588 N35589 Segment
X35589 N35589 N35590 Segment
X35590 N35590 N35591 Segment
X35591 N35591 N35592 Segment
X35592 N35592 N35593 Segment
X35593 N35593 N35594 Segment
X35594 N35594 N35595 Segment
X35595 N35595 N35596 Segment
X35596 N35596 N35597 Segment
X35597 N35597 N35598 Segment
X35598 N35598 N35599 Segment
X35599 N35599 N35600 Segment
X35600 N35600 N35601 Segment
X35601 N35601 N35602 Segment
X35602 N35602 N35603 Segment
X35603 N35603 N35604 Segment
X35604 N35604 N35605 Segment
X35605 N35605 N35606 Segment
X35606 N35606 N35607 Segment
X35607 N35607 N35608 Segment
X35608 N35608 N35609 Segment
X35609 N35609 N35610 Segment
X35610 N35610 N35611 Segment
X35611 N35611 N35612 Segment
X35612 N35612 N35613 Segment
X35613 N35613 N35614 Segment
X35614 N35614 N35615 Segment
X35615 N35615 N35616 Segment
X35616 N35616 N35617 Segment
X35617 N35617 N35618 Segment
X35618 N35618 N35619 Segment
X35619 N35619 N35620 Segment
X35620 N35620 N35621 Segment
X35621 N35621 N35622 Segment
X35622 N35622 N35623 Segment
X35623 N35623 N35624 Segment
X35624 N35624 N35625 Segment
X35625 N35625 N35626 Segment
X35626 N35626 N35627 Segment
X35627 N35627 N35628 Segment
X35628 N35628 N35629 Segment
X35629 N35629 N35630 Segment
X35630 N35630 N35631 Segment
X35631 N35631 N35632 Segment
X35632 N35632 N35633 Segment
X35633 N35633 N35634 Segment
X35634 N35634 N35635 Segment
X35635 N35635 N35636 Segment
X35636 N35636 N35637 Segment
X35637 N35637 N35638 Segment
X35638 N35638 N35639 Segment
X35639 N35639 N35640 Segment
X35640 N35640 N35641 Segment
X35641 N35641 N35642 Segment
X35642 N35642 N35643 Segment
X35643 N35643 N35644 Segment
X35644 N35644 N35645 Segment
X35645 N35645 N35646 Segment
X35646 N35646 N35647 Segment
X35647 N35647 N35648 Segment
X35648 N35648 N35649 Segment
X35649 N35649 N35650 Segment
X35650 N35650 N35651 Segment
X35651 N35651 N35652 Segment
X35652 N35652 N35653 Segment
X35653 N35653 N35654 Segment
X35654 N35654 N35655 Segment
X35655 N35655 N35656 Segment
X35656 N35656 N35657 Segment
X35657 N35657 N35658 Segment
X35658 N35658 N35659 Segment
X35659 N35659 N35660 Segment
X35660 N35660 N35661 Segment
X35661 N35661 N35662 Segment
X35662 N35662 N35663 Segment
X35663 N35663 N35664 Segment
X35664 N35664 N35665 Segment
X35665 N35665 N35666 Segment
X35666 N35666 N35667 Segment
X35667 N35667 N35668 Segment
X35668 N35668 N35669 Segment
X35669 N35669 N35670 Segment
X35670 N35670 N35671 Segment
X35671 N35671 N35672 Segment
X35672 N35672 N35673 Segment
X35673 N35673 N35674 Segment
X35674 N35674 N35675 Segment
X35675 N35675 N35676 Segment
X35676 N35676 N35677 Segment
X35677 N35677 N35678 Segment
X35678 N35678 N35679 Segment
X35679 N35679 N35680 Segment
X35680 N35680 N35681 Segment
X35681 N35681 N35682 Segment
X35682 N35682 N35683 Segment
X35683 N35683 N35684 Segment
X35684 N35684 N35685 Segment
X35685 N35685 N35686 Segment
X35686 N35686 N35687 Segment
X35687 N35687 N35688 Segment
X35688 N35688 N35689 Segment
X35689 N35689 N35690 Segment
X35690 N35690 N35691 Segment
X35691 N35691 N35692 Segment
X35692 N35692 N35693 Segment
X35693 N35693 N35694 Segment
X35694 N35694 N35695 Segment
X35695 N35695 N35696 Segment
X35696 N35696 N35697 Segment
X35697 N35697 N35698 Segment
X35698 N35698 N35699 Segment
X35699 N35699 N35700 Segment
X35700 N35700 N35701 Segment
X35701 N35701 N35702 Segment
X35702 N35702 N35703 Segment
X35703 N35703 N35704 Segment
X35704 N35704 N35705 Segment
X35705 N35705 N35706 Segment
X35706 N35706 N35707 Segment
X35707 N35707 N35708 Segment
X35708 N35708 N35709 Segment
X35709 N35709 N35710 Segment
X35710 N35710 N35711 Segment
X35711 N35711 N35712 Segment
X35712 N35712 N35713 Segment
X35713 N35713 N35714 Segment
X35714 N35714 N35715 Segment
X35715 N35715 N35716 Segment
X35716 N35716 N35717 Segment
X35717 N35717 N35718 Segment
X35718 N35718 N35719 Segment
X35719 N35719 N35720 Segment
X35720 N35720 N35721 Segment
X35721 N35721 N35722 Segment
X35722 N35722 N35723 Segment
X35723 N35723 N35724 Segment
X35724 N35724 N35725 Segment
X35725 N35725 N35726 Segment
X35726 N35726 N35727 Segment
X35727 N35727 N35728 Segment
X35728 N35728 N35729 Segment
X35729 N35729 N35730 Segment
X35730 N35730 N35731 Segment
X35731 N35731 N35732 Segment
X35732 N35732 N35733 Segment
X35733 N35733 N35734 Segment
X35734 N35734 N35735 Segment
X35735 N35735 N35736 Segment
X35736 N35736 N35737 Segment
X35737 N35737 N35738 Segment
X35738 N35738 N35739 Segment
X35739 N35739 N35740 Segment
X35740 N35740 N35741 Segment
X35741 N35741 N35742 Segment
X35742 N35742 N35743 Segment
X35743 N35743 N35744 Segment
X35744 N35744 N35745 Segment
X35745 N35745 N35746 Segment
X35746 N35746 N35747 Segment
X35747 N35747 N35748 Segment
X35748 N35748 N35749 Segment
X35749 N35749 N35750 Segment
X35750 N35750 N35751 Segment
X35751 N35751 N35752 Segment
X35752 N35752 N35753 Segment
X35753 N35753 N35754 Segment
X35754 N35754 N35755 Segment
X35755 N35755 N35756 Segment
X35756 N35756 N35757 Segment
X35757 N35757 N35758 Segment
X35758 N35758 N35759 Segment
X35759 N35759 N35760 Segment
X35760 N35760 N35761 Segment
X35761 N35761 N35762 Segment
X35762 N35762 N35763 Segment
X35763 N35763 N35764 Segment
X35764 N35764 N35765 Segment
X35765 N35765 N35766 Segment
X35766 N35766 N35767 Segment
X35767 N35767 N35768 Segment
X35768 N35768 N35769 Segment
X35769 N35769 N35770 Segment
X35770 N35770 N35771 Segment
X35771 N35771 N35772 Segment
X35772 N35772 N35773 Segment
X35773 N35773 N35774 Segment
X35774 N35774 N35775 Segment
X35775 N35775 N35776 Segment
X35776 N35776 N35777 Segment
X35777 N35777 N35778 Segment
X35778 N35778 N35779 Segment
X35779 N35779 N35780 Segment
X35780 N35780 N35781 Segment
X35781 N35781 N35782 Segment
X35782 N35782 N35783 Segment
X35783 N35783 N35784 Segment
X35784 N35784 N35785 Segment
X35785 N35785 N35786 Segment
X35786 N35786 N35787 Segment
X35787 N35787 N35788 Segment
X35788 N35788 N35789 Segment
X35789 N35789 N35790 Segment
X35790 N35790 N35791 Segment
X35791 N35791 N35792 Segment
X35792 N35792 N35793 Segment
X35793 N35793 N35794 Segment
X35794 N35794 N35795 Segment
X35795 N35795 N35796 Segment
X35796 N35796 N35797 Segment
X35797 N35797 N35798 Segment
X35798 N35798 N35799 Segment
X35799 N35799 N35800 Segment
X35800 N35800 N35801 Segment
X35801 N35801 N35802 Segment
X35802 N35802 N35803 Segment
X35803 N35803 N35804 Segment
X35804 N35804 N35805 Segment
X35805 N35805 N35806 Segment
X35806 N35806 N35807 Segment
X35807 N35807 N35808 Segment
X35808 N35808 N35809 Segment
X35809 N35809 N35810 Segment
X35810 N35810 N35811 Segment
X35811 N35811 N35812 Segment
X35812 N35812 N35813 Segment
X35813 N35813 N35814 Segment
X35814 N35814 N35815 Segment
X35815 N35815 N35816 Segment
X35816 N35816 N35817 Segment
X35817 N35817 N35818 Segment
X35818 N35818 N35819 Segment
X35819 N35819 N35820 Segment
X35820 N35820 N35821 Segment
X35821 N35821 N35822 Segment
X35822 N35822 N35823 Segment
X35823 N35823 N35824 Segment
X35824 N35824 N35825 Segment
X35825 N35825 N35826 Segment
X35826 N35826 N35827 Segment
X35827 N35827 N35828 Segment
X35828 N35828 N35829 Segment
X35829 N35829 N35830 Segment
X35830 N35830 N35831 Segment
X35831 N35831 N35832 Segment
X35832 N35832 N35833 Segment
X35833 N35833 N35834 Segment
X35834 N35834 N35835 Segment
X35835 N35835 N35836 Segment
X35836 N35836 N35837 Segment
X35837 N35837 N35838 Segment
X35838 N35838 N35839 Segment
X35839 N35839 N35840 Segment
X35840 N35840 N35841 Segment
X35841 N35841 N35842 Segment
X35842 N35842 N35843 Segment
X35843 N35843 N35844 Segment
X35844 N35844 N35845 Segment
X35845 N35845 N35846 Segment
X35846 N35846 N35847 Segment
X35847 N35847 N35848 Segment
X35848 N35848 N35849 Segment
X35849 N35849 N35850 Segment
X35850 N35850 N35851 Segment
X35851 N35851 N35852 Segment
X35852 N35852 N35853 Segment
X35853 N35853 N35854 Segment
X35854 N35854 N35855 Segment
X35855 N35855 N35856 Segment
X35856 N35856 N35857 Segment
X35857 N35857 N35858 Segment
X35858 N35858 N35859 Segment
X35859 N35859 N35860 Segment
X35860 N35860 N35861 Segment
X35861 N35861 N35862 Segment
X35862 N35862 N35863 Segment
X35863 N35863 N35864 Segment
X35864 N35864 N35865 Segment
X35865 N35865 N35866 Segment
X35866 N35866 N35867 Segment
X35867 N35867 N35868 Segment
X35868 N35868 N35869 Segment
X35869 N35869 N35870 Segment
X35870 N35870 N35871 Segment
X35871 N35871 N35872 Segment
X35872 N35872 N35873 Segment
X35873 N35873 N35874 Segment
X35874 N35874 N35875 Segment
X35875 N35875 N35876 Segment
X35876 N35876 N35877 Segment
X35877 N35877 N35878 Segment
X35878 N35878 N35879 Segment
X35879 N35879 N35880 Segment
X35880 N35880 N35881 Segment
X35881 N35881 N35882 Segment
X35882 N35882 N35883 Segment
X35883 N35883 N35884 Segment
X35884 N35884 N35885 Segment
X35885 N35885 N35886 Segment
X35886 N35886 N35887 Segment
X35887 N35887 N35888 Segment
X35888 N35888 N35889 Segment
X35889 N35889 N35890 Segment
X35890 N35890 N35891 Segment
X35891 N35891 N35892 Segment
X35892 N35892 N35893 Segment
X35893 N35893 N35894 Segment
X35894 N35894 N35895 Segment
X35895 N35895 N35896 Segment
X35896 N35896 N35897 Segment
X35897 N35897 N35898 Segment
X35898 N35898 N35899 Segment
X35899 N35899 N35900 Segment
X35900 N35900 N35901 Segment
X35901 N35901 N35902 Segment
X35902 N35902 N35903 Segment
X35903 N35903 N35904 Segment
X35904 N35904 N35905 Segment
X35905 N35905 N35906 Segment
X35906 N35906 N35907 Segment
X35907 N35907 N35908 Segment
X35908 N35908 N35909 Segment
X35909 N35909 N35910 Segment
X35910 N35910 N35911 Segment
X35911 N35911 N35912 Segment
X35912 N35912 N35913 Segment
X35913 N35913 N35914 Segment
X35914 N35914 N35915 Segment
X35915 N35915 N35916 Segment
X35916 N35916 N35917 Segment
X35917 N35917 N35918 Segment
X35918 N35918 N35919 Segment
X35919 N35919 N35920 Segment
X35920 N35920 N35921 Segment
X35921 N35921 N35922 Segment
X35922 N35922 N35923 Segment
X35923 N35923 N35924 Segment
X35924 N35924 N35925 Segment
X35925 N35925 N35926 Segment
X35926 N35926 N35927 Segment
X35927 N35927 N35928 Segment
X35928 N35928 N35929 Segment
X35929 N35929 N35930 Segment
X35930 N35930 N35931 Segment
X35931 N35931 N35932 Segment
X35932 N35932 N35933 Segment
X35933 N35933 N35934 Segment
X35934 N35934 N35935 Segment
X35935 N35935 N35936 Segment
X35936 N35936 N35937 Segment
X35937 N35937 N35938 Segment
X35938 N35938 N35939 Segment
X35939 N35939 N35940 Segment
X35940 N35940 N35941 Segment
X35941 N35941 N35942 Segment
X35942 N35942 N35943 Segment
X35943 N35943 N35944 Segment
X35944 N35944 N35945 Segment
X35945 N35945 N35946 Segment
X35946 N35946 N35947 Segment
X35947 N35947 N35948 Segment
X35948 N35948 N35949 Segment
X35949 N35949 N35950 Segment
X35950 N35950 N35951 Segment
X35951 N35951 N35952 Segment
X35952 N35952 N35953 Segment
X35953 N35953 N35954 Segment
X35954 N35954 N35955 Segment
X35955 N35955 N35956 Segment
X35956 N35956 N35957 Segment
X35957 N35957 N35958 Segment
X35958 N35958 N35959 Segment
X35959 N35959 N35960 Segment
X35960 N35960 N35961 Segment
X35961 N35961 N35962 Segment
X35962 N35962 N35963 Segment
X35963 N35963 N35964 Segment
X35964 N35964 N35965 Segment
X35965 N35965 N35966 Segment
X35966 N35966 N35967 Segment
X35967 N35967 N35968 Segment
X35968 N35968 N35969 Segment
X35969 N35969 N35970 Segment
X35970 N35970 N35971 Segment
X35971 N35971 N35972 Segment
X35972 N35972 N35973 Segment
X35973 N35973 N35974 Segment
X35974 N35974 N35975 Segment
X35975 N35975 N35976 Segment
X35976 N35976 N35977 Segment
X35977 N35977 N35978 Segment
X35978 N35978 N35979 Segment
X35979 N35979 N35980 Segment
X35980 N35980 N35981 Segment
X35981 N35981 N35982 Segment
X35982 N35982 N35983 Segment
X35983 N35983 N35984 Segment
X35984 N35984 N35985 Segment
X35985 N35985 N35986 Segment
X35986 N35986 N35987 Segment
X35987 N35987 N35988 Segment
X35988 N35988 N35989 Segment
X35989 N35989 N35990 Segment
X35990 N35990 N35991 Segment
X35991 N35991 N35992 Segment
X35992 N35992 N35993 Segment
X35993 N35993 N35994 Segment
X35994 N35994 N35995 Segment
X35995 N35995 N35996 Segment
X35996 N35996 N35997 Segment
X35997 N35997 N35998 Segment
X35998 N35998 N35999 Segment
X35999 N35999 N36000 Segment
X36000 N36000 N36001 Segment
X36001 N36001 N36002 Segment
X36002 N36002 N36003 Segment
X36003 N36003 N36004 Segment
X36004 N36004 N36005 Segment
X36005 N36005 N36006 Segment
X36006 N36006 N36007 Segment
X36007 N36007 N36008 Segment
X36008 N36008 N36009 Segment
X36009 N36009 N36010 Segment
X36010 N36010 N36011 Segment
X36011 N36011 N36012 Segment
X36012 N36012 N36013 Segment
X36013 N36013 N36014 Segment
X36014 N36014 N36015 Segment
X36015 N36015 N36016 Segment
X36016 N36016 N36017 Segment
X36017 N36017 N36018 Segment
X36018 N36018 N36019 Segment
X36019 N36019 N36020 Segment
X36020 N36020 N36021 Segment
X36021 N36021 N36022 Segment
X36022 N36022 N36023 Segment
X36023 N36023 N36024 Segment
X36024 N36024 N36025 Segment
X36025 N36025 N36026 Segment
X36026 N36026 N36027 Segment
X36027 N36027 N36028 Segment
X36028 N36028 N36029 Segment
X36029 N36029 N36030 Segment
X36030 N36030 N36031 Segment
X36031 N36031 N36032 Segment
X36032 N36032 N36033 Segment
X36033 N36033 N36034 Segment
X36034 N36034 N36035 Segment
X36035 N36035 N36036 Segment
X36036 N36036 N36037 Segment
X36037 N36037 N36038 Segment
X36038 N36038 N36039 Segment
X36039 N36039 N36040 Segment
X36040 N36040 N36041 Segment
X36041 N36041 N36042 Segment
X36042 N36042 N36043 Segment
X36043 N36043 N36044 Segment
X36044 N36044 N36045 Segment
X36045 N36045 N36046 Segment
X36046 N36046 N36047 Segment
X36047 N36047 N36048 Segment
X36048 N36048 N36049 Segment
X36049 N36049 N36050 Segment
X36050 N36050 N36051 Segment
X36051 N36051 N36052 Segment
X36052 N36052 N36053 Segment
X36053 N36053 N36054 Segment
X36054 N36054 N36055 Segment
X36055 N36055 N36056 Segment
X36056 N36056 N36057 Segment
X36057 N36057 N36058 Segment
X36058 N36058 N36059 Segment
X36059 N36059 N36060 Segment
X36060 N36060 N36061 Segment
X36061 N36061 N36062 Segment
X36062 N36062 N36063 Segment
X36063 N36063 N36064 Segment
X36064 N36064 N36065 Segment
X36065 N36065 N36066 Segment
X36066 N36066 N36067 Segment
X36067 N36067 N36068 Segment
X36068 N36068 N36069 Segment
X36069 N36069 N36070 Segment
X36070 N36070 N36071 Segment
X36071 N36071 N36072 Segment
X36072 N36072 N36073 Segment
X36073 N36073 N36074 Segment
X36074 N36074 N36075 Segment
X36075 N36075 N36076 Segment
X36076 N36076 N36077 Segment
X36077 N36077 N36078 Segment
X36078 N36078 N36079 Segment
X36079 N36079 N36080 Segment
X36080 N36080 N36081 Segment
X36081 N36081 N36082 Segment
X36082 N36082 N36083 Segment
X36083 N36083 N36084 Segment
X36084 N36084 N36085 Segment
X36085 N36085 N36086 Segment
X36086 N36086 N36087 Segment
X36087 N36087 N36088 Segment
X36088 N36088 N36089 Segment
X36089 N36089 N36090 Segment
X36090 N36090 N36091 Segment
X36091 N36091 N36092 Segment
X36092 N36092 N36093 Segment
X36093 N36093 N36094 Segment
X36094 N36094 N36095 Segment
X36095 N36095 N36096 Segment
X36096 N36096 N36097 Segment
X36097 N36097 N36098 Segment
X36098 N36098 N36099 Segment
X36099 N36099 N36100 Segment
X36100 N36100 N36101 Segment
X36101 N36101 N36102 Segment
X36102 N36102 N36103 Segment
X36103 N36103 N36104 Segment
X36104 N36104 N36105 Segment
X36105 N36105 N36106 Segment
X36106 N36106 N36107 Segment
X36107 N36107 N36108 Segment
X36108 N36108 N36109 Segment
X36109 N36109 N36110 Segment
X36110 N36110 N36111 Segment
X36111 N36111 N36112 Segment
X36112 N36112 N36113 Segment
X36113 N36113 N36114 Segment
X36114 N36114 N36115 Segment
X36115 N36115 N36116 Segment
X36116 N36116 N36117 Segment
X36117 N36117 N36118 Segment
X36118 N36118 N36119 Segment
X36119 N36119 N36120 Segment
X36120 N36120 N36121 Segment
X36121 N36121 N36122 Segment
X36122 N36122 N36123 Segment
X36123 N36123 N36124 Segment
X36124 N36124 N36125 Segment
X36125 N36125 N36126 Segment
X36126 N36126 N36127 Segment
X36127 N36127 N36128 Segment
X36128 N36128 N36129 Segment
X36129 N36129 N36130 Segment
X36130 N36130 N36131 Segment
X36131 N36131 N36132 Segment
X36132 N36132 N36133 Segment
X36133 N36133 N36134 Segment
X36134 N36134 N36135 Segment
X36135 N36135 N36136 Segment
X36136 N36136 N36137 Segment
X36137 N36137 N36138 Segment
X36138 N36138 N36139 Segment
X36139 N36139 N36140 Segment
X36140 N36140 N36141 Segment
X36141 N36141 N36142 Segment
X36142 N36142 N36143 Segment
X36143 N36143 N36144 Segment
X36144 N36144 N36145 Segment
X36145 N36145 N36146 Segment
X36146 N36146 N36147 Segment
X36147 N36147 N36148 Segment
X36148 N36148 N36149 Segment
X36149 N36149 N36150 Segment
X36150 N36150 N36151 Segment
X36151 N36151 N36152 Segment
X36152 N36152 N36153 Segment
X36153 N36153 N36154 Segment
X36154 N36154 N36155 Segment
X36155 N36155 N36156 Segment
X36156 N36156 N36157 Segment
X36157 N36157 N36158 Segment
X36158 N36158 N36159 Segment
X36159 N36159 N36160 Segment
X36160 N36160 N36161 Segment
X36161 N36161 N36162 Segment
X36162 N36162 N36163 Segment
X36163 N36163 N36164 Segment
X36164 N36164 N36165 Segment
X36165 N36165 N36166 Segment
X36166 N36166 N36167 Segment
X36167 N36167 N36168 Segment
X36168 N36168 N36169 Segment
X36169 N36169 N36170 Segment
X36170 N36170 N36171 Segment
X36171 N36171 N36172 Segment
X36172 N36172 N36173 Segment
X36173 N36173 N36174 Segment
X36174 N36174 N36175 Segment
X36175 N36175 N36176 Segment
X36176 N36176 N36177 Segment
X36177 N36177 N36178 Segment
X36178 N36178 N36179 Segment
X36179 N36179 N36180 Segment
X36180 N36180 N36181 Segment
X36181 N36181 N36182 Segment
X36182 N36182 N36183 Segment
X36183 N36183 N36184 Segment
X36184 N36184 N36185 Segment
X36185 N36185 N36186 Segment
X36186 N36186 N36187 Segment
X36187 N36187 N36188 Segment
X36188 N36188 N36189 Segment
X36189 N36189 N36190 Segment
X36190 N36190 N36191 Segment
X36191 N36191 N36192 Segment
X36192 N36192 N36193 Segment
X36193 N36193 N36194 Segment
X36194 N36194 N36195 Segment
X36195 N36195 N36196 Segment
X36196 N36196 N36197 Segment
X36197 N36197 N36198 Segment
X36198 N36198 N36199 Segment
X36199 N36199 N36200 Segment
X36200 N36200 N36201 Segment
X36201 N36201 N36202 Segment
X36202 N36202 N36203 Segment
X36203 N36203 N36204 Segment
X36204 N36204 N36205 Segment
X36205 N36205 N36206 Segment
X36206 N36206 N36207 Segment
X36207 N36207 N36208 Segment
X36208 N36208 N36209 Segment
X36209 N36209 N36210 Segment
X36210 N36210 N36211 Segment
X36211 N36211 N36212 Segment
X36212 N36212 N36213 Segment
X36213 N36213 N36214 Segment
X36214 N36214 N36215 Segment
X36215 N36215 N36216 Segment
X36216 N36216 N36217 Segment
X36217 N36217 N36218 Segment
X36218 N36218 N36219 Segment
X36219 N36219 N36220 Segment
X36220 N36220 N36221 Segment
X36221 N36221 N36222 Segment
X36222 N36222 N36223 Segment
X36223 N36223 N36224 Segment
X36224 N36224 N36225 Segment
X36225 N36225 N36226 Segment
X36226 N36226 N36227 Segment
X36227 N36227 N36228 Segment
X36228 N36228 N36229 Segment
X36229 N36229 N36230 Segment
X36230 N36230 N36231 Segment
X36231 N36231 N36232 Segment
X36232 N36232 N36233 Segment
X36233 N36233 N36234 Segment
X36234 N36234 N36235 Segment
X36235 N36235 N36236 Segment
X36236 N36236 N36237 Segment
X36237 N36237 N36238 Segment
X36238 N36238 N36239 Segment
X36239 N36239 N36240 Segment
X36240 N36240 N36241 Segment
X36241 N36241 N36242 Segment
X36242 N36242 N36243 Segment
X36243 N36243 N36244 Segment
X36244 N36244 N36245 Segment
X36245 N36245 N36246 Segment
X36246 N36246 N36247 Segment
X36247 N36247 N36248 Segment
X36248 N36248 N36249 Segment
X36249 N36249 N36250 Segment
X36250 N36250 N36251 Segment
X36251 N36251 N36252 Segment
X36252 N36252 N36253 Segment
X36253 N36253 N36254 Segment
X36254 N36254 N36255 Segment
X36255 N36255 N36256 Segment
X36256 N36256 N36257 Segment
X36257 N36257 N36258 Segment
X36258 N36258 N36259 Segment
X36259 N36259 N36260 Segment
X36260 N36260 N36261 Segment
X36261 N36261 N36262 Segment
X36262 N36262 N36263 Segment
X36263 N36263 N36264 Segment
X36264 N36264 N36265 Segment
X36265 N36265 N36266 Segment
X36266 N36266 N36267 Segment
X36267 N36267 N36268 Segment
X36268 N36268 N36269 Segment
X36269 N36269 N36270 Segment
X36270 N36270 N36271 Segment
X36271 N36271 N36272 Segment
X36272 N36272 N36273 Segment
X36273 N36273 N36274 Segment
X36274 N36274 N36275 Segment
X36275 N36275 N36276 Segment
X36276 N36276 N36277 Segment
X36277 N36277 N36278 Segment
X36278 N36278 N36279 Segment
X36279 N36279 N36280 Segment
X36280 N36280 N36281 Segment
X36281 N36281 N36282 Segment
X36282 N36282 N36283 Segment
X36283 N36283 N36284 Segment
X36284 N36284 N36285 Segment
X36285 N36285 N36286 Segment
X36286 N36286 N36287 Segment
X36287 N36287 N36288 Segment
X36288 N36288 N36289 Segment
X36289 N36289 N36290 Segment
X36290 N36290 N36291 Segment
X36291 N36291 N36292 Segment
X36292 N36292 N36293 Segment
X36293 N36293 N36294 Segment
X36294 N36294 N36295 Segment
X36295 N36295 N36296 Segment
X36296 N36296 N36297 Segment
X36297 N36297 N36298 Segment
X36298 N36298 N36299 Segment
X36299 N36299 N36300 Segment
X36300 N36300 N36301 Segment
X36301 N36301 N36302 Segment
X36302 N36302 N36303 Segment
X36303 N36303 N36304 Segment
X36304 N36304 N36305 Segment
X36305 N36305 N36306 Segment
X36306 N36306 N36307 Segment
X36307 N36307 N36308 Segment
X36308 N36308 N36309 Segment
X36309 N36309 N36310 Segment
X36310 N36310 N36311 Segment
X36311 N36311 N36312 Segment
X36312 N36312 N36313 Segment
X36313 N36313 N36314 Segment
X36314 N36314 N36315 Segment
X36315 N36315 N36316 Segment
X36316 N36316 N36317 Segment
X36317 N36317 N36318 Segment
X36318 N36318 N36319 Segment
X36319 N36319 N36320 Segment
X36320 N36320 N36321 Segment
X36321 N36321 N36322 Segment
X36322 N36322 N36323 Segment
X36323 N36323 N36324 Segment
X36324 N36324 N36325 Segment
X36325 N36325 N36326 Segment
X36326 N36326 N36327 Segment
X36327 N36327 N36328 Segment
X36328 N36328 N36329 Segment
X36329 N36329 N36330 Segment
X36330 N36330 N36331 Segment
X36331 N36331 N36332 Segment
X36332 N36332 N36333 Segment
X36333 N36333 N36334 Segment
X36334 N36334 N36335 Segment
X36335 N36335 N36336 Segment
X36336 N36336 N36337 Segment
X36337 N36337 N36338 Segment
X36338 N36338 N36339 Segment
X36339 N36339 N36340 Segment
X36340 N36340 N36341 Segment
X36341 N36341 N36342 Segment
X36342 N36342 N36343 Segment
X36343 N36343 N36344 Segment
X36344 N36344 N36345 Segment
X36345 N36345 N36346 Segment
X36346 N36346 N36347 Segment
X36347 N36347 N36348 Segment
X36348 N36348 N36349 Segment
X36349 N36349 N36350 Segment
X36350 N36350 N36351 Segment
X36351 N36351 N36352 Segment
X36352 N36352 N36353 Segment
X36353 N36353 N36354 Segment
X36354 N36354 N36355 Segment
X36355 N36355 N36356 Segment
X36356 N36356 N36357 Segment
X36357 N36357 N36358 Segment
X36358 N36358 N36359 Segment
X36359 N36359 N36360 Segment
X36360 N36360 N36361 Segment
X36361 N36361 N36362 Segment
X36362 N36362 N36363 Segment
X36363 N36363 N36364 Segment
X36364 N36364 N36365 Segment
X36365 N36365 N36366 Segment
X36366 N36366 N36367 Segment
X36367 N36367 N36368 Segment
X36368 N36368 N36369 Segment
X36369 N36369 N36370 Segment
X36370 N36370 N36371 Segment
X36371 N36371 N36372 Segment
X36372 N36372 N36373 Segment
X36373 N36373 N36374 Segment
X36374 N36374 N36375 Segment
X36375 N36375 N36376 Segment
X36376 N36376 N36377 Segment
X36377 N36377 N36378 Segment
X36378 N36378 N36379 Segment
X36379 N36379 N36380 Segment
X36380 N36380 N36381 Segment
X36381 N36381 N36382 Segment
X36382 N36382 N36383 Segment
X36383 N36383 N36384 Segment
X36384 N36384 N36385 Segment
X36385 N36385 N36386 Segment
X36386 N36386 N36387 Segment
X36387 N36387 N36388 Segment
X36388 N36388 N36389 Segment
X36389 N36389 N36390 Segment
X36390 N36390 N36391 Segment
X36391 N36391 N36392 Segment
X36392 N36392 N36393 Segment
X36393 N36393 N36394 Segment
X36394 N36394 N36395 Segment
X36395 N36395 N36396 Segment
X36396 N36396 N36397 Segment
X36397 N36397 N36398 Segment
X36398 N36398 N36399 Segment
X36399 N36399 N36400 Segment
X36400 N36400 N36401 Segment
X36401 N36401 N36402 Segment
X36402 N36402 N36403 Segment
X36403 N36403 N36404 Segment
X36404 N36404 N36405 Segment
X36405 N36405 N36406 Segment
X36406 N36406 N36407 Segment
X36407 N36407 N36408 Segment
X36408 N36408 N36409 Segment
X36409 N36409 N36410 Segment
X36410 N36410 N36411 Segment
X36411 N36411 N36412 Segment
X36412 N36412 N36413 Segment
X36413 N36413 N36414 Segment
X36414 N36414 N36415 Segment
X36415 N36415 N36416 Segment
X36416 N36416 N36417 Segment
X36417 N36417 N36418 Segment
X36418 N36418 N36419 Segment
X36419 N36419 N36420 Segment
X36420 N36420 N36421 Segment
X36421 N36421 N36422 Segment
X36422 N36422 N36423 Segment
X36423 N36423 N36424 Segment
X36424 N36424 N36425 Segment
X36425 N36425 N36426 Segment
X36426 N36426 N36427 Segment
X36427 N36427 N36428 Segment
X36428 N36428 N36429 Segment
X36429 N36429 N36430 Segment
X36430 N36430 N36431 Segment
X36431 N36431 N36432 Segment
X36432 N36432 N36433 Segment
X36433 N36433 N36434 Segment
X36434 N36434 N36435 Segment
X36435 N36435 N36436 Segment
X36436 N36436 N36437 Segment
X36437 N36437 N36438 Segment
X36438 N36438 N36439 Segment
X36439 N36439 N36440 Segment
X36440 N36440 N36441 Segment
X36441 N36441 N36442 Segment
X36442 N36442 N36443 Segment
X36443 N36443 N36444 Segment
X36444 N36444 N36445 Segment
X36445 N36445 N36446 Segment
X36446 N36446 N36447 Segment
X36447 N36447 N36448 Segment
X36448 N36448 N36449 Segment
X36449 N36449 N36450 Segment
X36450 N36450 N36451 Segment
X36451 N36451 N36452 Segment
X36452 N36452 N36453 Segment
X36453 N36453 N36454 Segment
X36454 N36454 N36455 Segment
X36455 N36455 N36456 Segment
X36456 N36456 N36457 Segment
X36457 N36457 N36458 Segment
X36458 N36458 N36459 Segment
X36459 N36459 N36460 Segment
X36460 N36460 N36461 Segment
X36461 N36461 N36462 Segment
X36462 N36462 N36463 Segment
X36463 N36463 N36464 Segment
X36464 N36464 N36465 Segment
X36465 N36465 N36466 Segment
X36466 N36466 N36467 Segment
X36467 N36467 N36468 Segment
X36468 N36468 N36469 Segment
X36469 N36469 N36470 Segment
X36470 N36470 N36471 Segment
X36471 N36471 N36472 Segment
X36472 N36472 N36473 Segment
X36473 N36473 N36474 Segment
X36474 N36474 N36475 Segment
X36475 N36475 N36476 Segment
X36476 N36476 N36477 Segment
X36477 N36477 N36478 Segment
X36478 N36478 N36479 Segment
X36479 N36479 N36480 Segment
X36480 N36480 N36481 Segment
X36481 N36481 N36482 Segment
X36482 N36482 N36483 Segment
X36483 N36483 N36484 Segment
X36484 N36484 N36485 Segment
X36485 N36485 N36486 Segment
X36486 N36486 N36487 Segment
X36487 N36487 N36488 Segment
X36488 N36488 N36489 Segment
X36489 N36489 N36490 Segment
X36490 N36490 N36491 Segment
X36491 N36491 N36492 Segment
X36492 N36492 N36493 Segment
X36493 N36493 N36494 Segment
X36494 N36494 N36495 Segment
X36495 N36495 N36496 Segment
X36496 N36496 N36497 Segment
X36497 N36497 N36498 Segment
X36498 N36498 N36499 Segment
X36499 N36499 N36500 Segment
X36500 N36500 N36501 Segment
X36501 N36501 N36502 Segment
X36502 N36502 N36503 Segment
X36503 N36503 N36504 Segment
X36504 N36504 N36505 Segment
X36505 N36505 N36506 Segment
X36506 N36506 N36507 Segment
X36507 N36507 N36508 Segment
X36508 N36508 N36509 Segment
X36509 N36509 N36510 Segment
X36510 N36510 N36511 Segment
X36511 N36511 N36512 Segment
X36512 N36512 N36513 Segment
X36513 N36513 N36514 Segment
X36514 N36514 N36515 Segment
X36515 N36515 N36516 Segment
X36516 N36516 N36517 Segment
X36517 N36517 N36518 Segment
X36518 N36518 N36519 Segment
X36519 N36519 N36520 Segment
X36520 N36520 N36521 Segment
X36521 N36521 N36522 Segment
X36522 N36522 N36523 Segment
X36523 N36523 N36524 Segment
X36524 N36524 N36525 Segment
X36525 N36525 N36526 Segment
X36526 N36526 N36527 Segment
X36527 N36527 N36528 Segment
X36528 N36528 N36529 Segment
X36529 N36529 N36530 Segment
X36530 N36530 N36531 Segment
X36531 N36531 N36532 Segment
X36532 N36532 N36533 Segment
X36533 N36533 N36534 Segment
X36534 N36534 N36535 Segment
X36535 N36535 N36536 Segment
X36536 N36536 N36537 Segment
X36537 N36537 N36538 Segment
X36538 N36538 N36539 Segment
X36539 N36539 N36540 Segment
X36540 N36540 N36541 Segment
X36541 N36541 N36542 Segment
X36542 N36542 N36543 Segment
X36543 N36543 N36544 Segment
X36544 N36544 N36545 Segment
X36545 N36545 N36546 Segment
X36546 N36546 N36547 Segment
X36547 N36547 N36548 Segment
X36548 N36548 N36549 Segment
X36549 N36549 N36550 Segment
X36550 N36550 N36551 Segment
X36551 N36551 N36552 Segment
X36552 N36552 N36553 Segment
X36553 N36553 N36554 Segment
X36554 N36554 N36555 Segment
X36555 N36555 N36556 Segment
X36556 N36556 N36557 Segment
X36557 N36557 N36558 Segment
X36558 N36558 N36559 Segment
X36559 N36559 N36560 Segment
X36560 N36560 N36561 Segment
X36561 N36561 N36562 Segment
X36562 N36562 N36563 Segment
X36563 N36563 N36564 Segment
X36564 N36564 N36565 Segment
X36565 N36565 N36566 Segment
X36566 N36566 N36567 Segment
X36567 N36567 N36568 Segment
X36568 N36568 N36569 Segment
X36569 N36569 N36570 Segment
X36570 N36570 N36571 Segment
X36571 N36571 N36572 Segment
X36572 N36572 N36573 Segment
X36573 N36573 N36574 Segment
X36574 N36574 N36575 Segment
X36575 N36575 N36576 Segment
X36576 N36576 N36577 Segment
X36577 N36577 N36578 Segment
X36578 N36578 N36579 Segment
X36579 N36579 N36580 Segment
X36580 N36580 N36581 Segment
X36581 N36581 N36582 Segment
X36582 N36582 N36583 Segment
X36583 N36583 N36584 Segment
X36584 N36584 N36585 Segment
X36585 N36585 N36586 Segment
X36586 N36586 N36587 Segment
X36587 N36587 N36588 Segment
X36588 N36588 N36589 Segment
X36589 N36589 N36590 Segment
X36590 N36590 N36591 Segment
X36591 N36591 N36592 Segment
X36592 N36592 N36593 Segment
X36593 N36593 N36594 Segment
X36594 N36594 N36595 Segment
X36595 N36595 N36596 Segment
X36596 N36596 N36597 Segment
X36597 N36597 N36598 Segment
X36598 N36598 N36599 Segment
X36599 N36599 N36600 Segment
X36600 N36600 N36601 Segment
X36601 N36601 N36602 Segment
X36602 N36602 N36603 Segment
X36603 N36603 N36604 Segment
X36604 N36604 N36605 Segment
X36605 N36605 N36606 Segment
X36606 N36606 N36607 Segment
X36607 N36607 N36608 Segment
X36608 N36608 N36609 Segment
X36609 N36609 N36610 Segment
X36610 N36610 N36611 Segment
X36611 N36611 N36612 Segment
X36612 N36612 N36613 Segment
X36613 N36613 N36614 Segment
X36614 N36614 N36615 Segment
X36615 N36615 N36616 Segment
X36616 N36616 N36617 Segment
X36617 N36617 N36618 Segment
X36618 N36618 N36619 Segment
X36619 N36619 N36620 Segment
X36620 N36620 N36621 Segment
X36621 N36621 N36622 Segment
X36622 N36622 N36623 Segment
X36623 N36623 N36624 Segment
X36624 N36624 N36625 Segment
X36625 N36625 N36626 Segment
X36626 N36626 N36627 Segment
X36627 N36627 N36628 Segment
X36628 N36628 N36629 Segment
X36629 N36629 N36630 Segment
X36630 N36630 N36631 Segment
X36631 N36631 N36632 Segment
X36632 N36632 N36633 Segment
X36633 N36633 N36634 Segment
X36634 N36634 N36635 Segment
X36635 N36635 N36636 Segment
X36636 N36636 N36637 Segment
X36637 N36637 N36638 Segment
X36638 N36638 N36639 Segment
X36639 N36639 N36640 Segment
X36640 N36640 N36641 Segment
X36641 N36641 N36642 Segment
X36642 N36642 N36643 Segment
X36643 N36643 N36644 Segment
X36644 N36644 N36645 Segment
X36645 N36645 N36646 Segment
X36646 N36646 N36647 Segment
X36647 N36647 N36648 Segment
X36648 N36648 N36649 Segment
X36649 N36649 N36650 Segment
X36650 N36650 N36651 Segment
X36651 N36651 N36652 Segment
X36652 N36652 N36653 Segment
X36653 N36653 N36654 Segment
X36654 N36654 N36655 Segment
X36655 N36655 N36656 Segment
X36656 N36656 N36657 Segment
X36657 N36657 N36658 Segment
X36658 N36658 N36659 Segment
X36659 N36659 N36660 Segment
X36660 N36660 N36661 Segment
X36661 N36661 N36662 Segment
X36662 N36662 N36663 Segment
X36663 N36663 N36664 Segment
X36664 N36664 N36665 Segment
X36665 N36665 N36666 Segment
X36666 N36666 N36667 Segment
X36667 N36667 N36668 Segment
X36668 N36668 N36669 Segment
X36669 N36669 N36670 Segment
X36670 N36670 N36671 Segment
X36671 N36671 N36672 Segment
X36672 N36672 N36673 Segment
X36673 N36673 N36674 Segment
X36674 N36674 N36675 Segment
X36675 N36675 N36676 Segment
X36676 N36676 N36677 Segment
X36677 N36677 N36678 Segment
X36678 N36678 N36679 Segment
X36679 N36679 N36680 Segment
X36680 N36680 N36681 Segment
X36681 N36681 N36682 Segment
X36682 N36682 N36683 Segment
X36683 N36683 N36684 Segment
X36684 N36684 N36685 Segment
X36685 N36685 N36686 Segment
X36686 N36686 N36687 Segment
X36687 N36687 N36688 Segment
X36688 N36688 N36689 Segment
X36689 N36689 N36690 Segment
X36690 N36690 N36691 Segment
X36691 N36691 N36692 Segment
X36692 N36692 N36693 Segment
X36693 N36693 N36694 Segment
X36694 N36694 N36695 Segment
X36695 N36695 N36696 Segment
X36696 N36696 N36697 Segment
X36697 N36697 N36698 Segment
X36698 N36698 N36699 Segment
X36699 N36699 N36700 Segment
X36700 N36700 N36701 Segment
X36701 N36701 N36702 Segment
X36702 N36702 N36703 Segment
X36703 N36703 N36704 Segment
X36704 N36704 N36705 Segment
X36705 N36705 N36706 Segment
X36706 N36706 N36707 Segment
X36707 N36707 N36708 Segment
X36708 N36708 N36709 Segment
X36709 N36709 N36710 Segment
X36710 N36710 N36711 Segment
X36711 N36711 N36712 Segment
X36712 N36712 N36713 Segment
X36713 N36713 N36714 Segment
X36714 N36714 N36715 Segment
X36715 N36715 N36716 Segment
X36716 N36716 N36717 Segment
X36717 N36717 N36718 Segment
X36718 N36718 N36719 Segment
X36719 N36719 N36720 Segment
X36720 N36720 N36721 Segment
X36721 N36721 N36722 Segment
X36722 N36722 N36723 Segment
X36723 N36723 N36724 Segment
X36724 N36724 N36725 Segment
X36725 N36725 N36726 Segment
X36726 N36726 N36727 Segment
X36727 N36727 N36728 Segment
X36728 N36728 N36729 Segment
X36729 N36729 N36730 Segment
X36730 N36730 N36731 Segment
X36731 N36731 N36732 Segment
X36732 N36732 N36733 Segment
X36733 N36733 N36734 Segment
X36734 N36734 N36735 Segment
X36735 N36735 N36736 Segment
X36736 N36736 N36737 Segment
X36737 N36737 N36738 Segment
X36738 N36738 N36739 Segment
X36739 N36739 N36740 Segment
X36740 N36740 N36741 Segment
X36741 N36741 N36742 Segment
X36742 N36742 N36743 Segment
X36743 N36743 N36744 Segment
X36744 N36744 N36745 Segment
X36745 N36745 N36746 Segment
X36746 N36746 N36747 Segment
X36747 N36747 N36748 Segment
X36748 N36748 N36749 Segment
X36749 N36749 N36750 Segment
X36750 N36750 N36751 Segment
X36751 N36751 N36752 Segment
X36752 N36752 N36753 Segment
X36753 N36753 N36754 Segment
X36754 N36754 N36755 Segment
X36755 N36755 N36756 Segment
X36756 N36756 N36757 Segment
X36757 N36757 N36758 Segment
X36758 N36758 N36759 Segment
X36759 N36759 N36760 Segment
X36760 N36760 N36761 Segment
X36761 N36761 N36762 Segment
X36762 N36762 N36763 Segment
X36763 N36763 N36764 Segment
X36764 N36764 N36765 Segment
X36765 N36765 N36766 Segment
X36766 N36766 N36767 Segment
X36767 N36767 N36768 Segment
X36768 N36768 N36769 Segment
X36769 N36769 N36770 Segment
X36770 N36770 N36771 Segment
X36771 N36771 N36772 Segment
X36772 N36772 N36773 Segment
X36773 N36773 N36774 Segment
X36774 N36774 N36775 Segment
X36775 N36775 N36776 Segment
X36776 N36776 N36777 Segment
X36777 N36777 N36778 Segment
X36778 N36778 N36779 Segment
X36779 N36779 N36780 Segment
X36780 N36780 N36781 Segment
X36781 N36781 N36782 Segment
X36782 N36782 N36783 Segment
X36783 N36783 N36784 Segment
X36784 N36784 N36785 Segment
X36785 N36785 N36786 Segment
X36786 N36786 N36787 Segment
X36787 N36787 N36788 Segment
X36788 N36788 N36789 Segment
X36789 N36789 N36790 Segment
X36790 N36790 N36791 Segment
X36791 N36791 N36792 Segment
X36792 N36792 N36793 Segment
X36793 N36793 N36794 Segment
X36794 N36794 N36795 Segment
X36795 N36795 N36796 Segment
X36796 N36796 N36797 Segment
X36797 N36797 N36798 Segment
X36798 N36798 N36799 Segment
X36799 N36799 N36800 Segment
X36800 N36800 N36801 Segment
X36801 N36801 N36802 Segment
X36802 N36802 N36803 Segment
X36803 N36803 N36804 Segment
X36804 N36804 N36805 Segment
X36805 N36805 N36806 Segment
X36806 N36806 N36807 Segment
X36807 N36807 N36808 Segment
X36808 N36808 N36809 Segment
X36809 N36809 N36810 Segment
X36810 N36810 N36811 Segment
X36811 N36811 N36812 Segment
X36812 N36812 N36813 Segment
X36813 N36813 N36814 Segment
X36814 N36814 N36815 Segment
X36815 N36815 N36816 Segment
X36816 N36816 N36817 Segment
X36817 N36817 N36818 Segment
X36818 N36818 N36819 Segment
X36819 N36819 N36820 Segment
X36820 N36820 N36821 Segment
X36821 N36821 N36822 Segment
X36822 N36822 N36823 Segment
X36823 N36823 N36824 Segment
X36824 N36824 N36825 Segment
X36825 N36825 N36826 Segment
X36826 N36826 N36827 Segment
X36827 N36827 N36828 Segment
X36828 N36828 N36829 Segment
X36829 N36829 N36830 Segment
X36830 N36830 N36831 Segment
X36831 N36831 N36832 Segment
X36832 N36832 N36833 Segment
X36833 N36833 N36834 Segment
X36834 N36834 N36835 Segment
X36835 N36835 N36836 Segment
X36836 N36836 N36837 Segment
X36837 N36837 N36838 Segment
X36838 N36838 N36839 Segment
X36839 N36839 N36840 Segment
X36840 N36840 N36841 Segment
X36841 N36841 N36842 Segment
X36842 N36842 N36843 Segment
X36843 N36843 N36844 Segment
X36844 N36844 N36845 Segment
X36845 N36845 N36846 Segment
X36846 N36846 N36847 Segment
X36847 N36847 N36848 Segment
X36848 N36848 N36849 Segment
X36849 N36849 N36850 Segment
X36850 N36850 N36851 Segment
X36851 N36851 N36852 Segment
X36852 N36852 N36853 Segment
X36853 N36853 N36854 Segment
X36854 N36854 N36855 Segment
X36855 N36855 N36856 Segment
X36856 N36856 N36857 Segment
X36857 N36857 N36858 Segment
X36858 N36858 N36859 Segment
X36859 N36859 N36860 Segment
X36860 N36860 N36861 Segment
X36861 N36861 N36862 Segment
X36862 N36862 N36863 Segment
X36863 N36863 N36864 Segment
X36864 N36864 N36865 Segment
X36865 N36865 N36866 Segment
X36866 N36866 N36867 Segment
X36867 N36867 N36868 Segment
X36868 N36868 N36869 Segment
X36869 N36869 N36870 Segment
X36870 N36870 N36871 Segment
X36871 N36871 N36872 Segment
X36872 N36872 N36873 Segment
X36873 N36873 N36874 Segment
X36874 N36874 N36875 Segment
X36875 N36875 N36876 Segment
X36876 N36876 N36877 Segment
X36877 N36877 N36878 Segment
X36878 N36878 N36879 Segment
X36879 N36879 N36880 Segment
X36880 N36880 N36881 Segment
X36881 N36881 N36882 Segment
X36882 N36882 N36883 Segment
X36883 N36883 N36884 Segment
X36884 N36884 N36885 Segment
X36885 N36885 N36886 Segment
X36886 N36886 N36887 Segment
X36887 N36887 N36888 Segment
X36888 N36888 N36889 Segment
X36889 N36889 N36890 Segment
X36890 N36890 N36891 Segment
X36891 N36891 N36892 Segment
X36892 N36892 N36893 Segment
X36893 N36893 N36894 Segment
X36894 N36894 N36895 Segment
X36895 N36895 N36896 Segment
X36896 N36896 N36897 Segment
X36897 N36897 N36898 Segment
X36898 N36898 N36899 Segment
X36899 N36899 N36900 Segment
X36900 N36900 N36901 Segment
X36901 N36901 N36902 Segment
X36902 N36902 N36903 Segment
X36903 N36903 N36904 Segment
X36904 N36904 N36905 Segment
X36905 N36905 N36906 Segment
X36906 N36906 N36907 Segment
X36907 N36907 N36908 Segment
X36908 N36908 N36909 Segment
X36909 N36909 N36910 Segment
X36910 N36910 N36911 Segment
X36911 N36911 N36912 Segment
X36912 N36912 N36913 Segment
X36913 N36913 N36914 Segment
X36914 N36914 N36915 Segment
X36915 N36915 N36916 Segment
X36916 N36916 N36917 Segment
X36917 N36917 N36918 Segment
X36918 N36918 N36919 Segment
X36919 N36919 N36920 Segment
X36920 N36920 N36921 Segment
X36921 N36921 N36922 Segment
X36922 N36922 N36923 Segment
X36923 N36923 N36924 Segment
X36924 N36924 N36925 Segment
X36925 N36925 N36926 Segment
X36926 N36926 N36927 Segment
X36927 N36927 N36928 Segment
X36928 N36928 N36929 Segment
X36929 N36929 N36930 Segment
X36930 N36930 N36931 Segment
X36931 N36931 N36932 Segment
X36932 N36932 N36933 Segment
X36933 N36933 N36934 Segment
X36934 N36934 N36935 Segment
X36935 N36935 N36936 Segment
X36936 N36936 N36937 Segment
X36937 N36937 N36938 Segment
X36938 N36938 N36939 Segment
X36939 N36939 N36940 Segment
X36940 N36940 N36941 Segment
X36941 N36941 N36942 Segment
X36942 N36942 N36943 Segment
X36943 N36943 N36944 Segment
X36944 N36944 N36945 Segment
X36945 N36945 N36946 Segment
X36946 N36946 N36947 Segment
X36947 N36947 N36948 Segment
X36948 N36948 N36949 Segment
X36949 N36949 N36950 Segment
X36950 N36950 N36951 Segment
X36951 N36951 N36952 Segment
X36952 N36952 N36953 Segment
X36953 N36953 N36954 Segment
X36954 N36954 N36955 Segment
X36955 N36955 N36956 Segment
X36956 N36956 N36957 Segment
X36957 N36957 N36958 Segment
X36958 N36958 N36959 Segment
X36959 N36959 N36960 Segment
X36960 N36960 N36961 Segment
X36961 N36961 N36962 Segment
X36962 N36962 N36963 Segment
X36963 N36963 N36964 Segment
X36964 N36964 N36965 Segment
X36965 N36965 N36966 Segment
X36966 N36966 N36967 Segment
X36967 N36967 N36968 Segment
X36968 N36968 N36969 Segment
X36969 N36969 N36970 Segment
X36970 N36970 N36971 Segment
X36971 N36971 N36972 Segment
X36972 N36972 N36973 Segment
X36973 N36973 N36974 Segment
X36974 N36974 N36975 Segment
X36975 N36975 N36976 Segment
X36976 N36976 N36977 Segment
X36977 N36977 N36978 Segment
X36978 N36978 N36979 Segment
X36979 N36979 N36980 Segment
X36980 N36980 N36981 Segment
X36981 N36981 N36982 Segment
X36982 N36982 N36983 Segment
X36983 N36983 N36984 Segment
X36984 N36984 N36985 Segment
X36985 N36985 N36986 Segment
X36986 N36986 N36987 Segment
X36987 N36987 N36988 Segment
X36988 N36988 N36989 Segment
X36989 N36989 N36990 Segment
X36990 N36990 N36991 Segment
X36991 N36991 N36992 Segment
X36992 N36992 N36993 Segment
X36993 N36993 N36994 Segment
X36994 N36994 N36995 Segment
X36995 N36995 N36996 Segment
X36996 N36996 N36997 Segment
X36997 N36997 N36998 Segment
X36998 N36998 N36999 Segment
X36999 N36999 N37000 Segment
X37000 N37000 N37001 Segment
X37001 N37001 N37002 Segment
X37002 N37002 N37003 Segment
X37003 N37003 N37004 Segment
X37004 N37004 N37005 Segment
X37005 N37005 N37006 Segment
X37006 N37006 N37007 Segment
X37007 N37007 N37008 Segment
X37008 N37008 N37009 Segment
X37009 N37009 N37010 Segment
X37010 N37010 N37011 Segment
X37011 N37011 N37012 Segment
X37012 N37012 N37013 Segment
X37013 N37013 N37014 Segment
X37014 N37014 N37015 Segment
X37015 N37015 N37016 Segment
X37016 N37016 N37017 Segment
X37017 N37017 N37018 Segment
X37018 N37018 N37019 Segment
X37019 N37019 N37020 Segment
X37020 N37020 N37021 Segment
X37021 N37021 N37022 Segment
X37022 N37022 N37023 Segment
X37023 N37023 N37024 Segment
X37024 N37024 N37025 Segment
X37025 N37025 N37026 Segment
X37026 N37026 N37027 Segment
X37027 N37027 N37028 Segment
X37028 N37028 N37029 Segment
X37029 N37029 N37030 Segment
X37030 N37030 N37031 Segment
X37031 N37031 N37032 Segment
X37032 N37032 N37033 Segment
X37033 N37033 N37034 Segment
X37034 N37034 N37035 Segment
X37035 N37035 N37036 Segment
X37036 N37036 N37037 Segment
X37037 N37037 N37038 Segment
X37038 N37038 N37039 Segment
X37039 N37039 N37040 Segment
X37040 N37040 N37041 Segment
X37041 N37041 N37042 Segment
X37042 N37042 N37043 Segment
X37043 N37043 N37044 Segment
X37044 N37044 N37045 Segment
X37045 N37045 N37046 Segment
X37046 N37046 N37047 Segment
X37047 N37047 N37048 Segment
X37048 N37048 N37049 Segment
X37049 N37049 N37050 Segment
X37050 N37050 N37051 Segment
X37051 N37051 N37052 Segment
X37052 N37052 N37053 Segment
X37053 N37053 N37054 Segment
X37054 N37054 N37055 Segment
X37055 N37055 N37056 Segment
X37056 N37056 N37057 Segment
X37057 N37057 N37058 Segment
X37058 N37058 N37059 Segment
X37059 N37059 N37060 Segment
X37060 N37060 N37061 Segment
X37061 N37061 N37062 Segment
X37062 N37062 N37063 Segment
X37063 N37063 N37064 Segment
X37064 N37064 N37065 Segment
X37065 N37065 N37066 Segment
X37066 N37066 N37067 Segment
X37067 N37067 N37068 Segment
X37068 N37068 N37069 Segment
X37069 N37069 N37070 Segment
X37070 N37070 N37071 Segment
X37071 N37071 N37072 Segment
X37072 N37072 N37073 Segment
X37073 N37073 N37074 Segment
X37074 N37074 N37075 Segment
X37075 N37075 N37076 Segment
X37076 N37076 N37077 Segment
X37077 N37077 N37078 Segment
X37078 N37078 N37079 Segment
X37079 N37079 N37080 Segment
X37080 N37080 N37081 Segment
X37081 N37081 N37082 Segment
X37082 N37082 N37083 Segment
X37083 N37083 N37084 Segment
X37084 N37084 N37085 Segment
X37085 N37085 N37086 Segment
X37086 N37086 N37087 Segment
X37087 N37087 N37088 Segment
X37088 N37088 N37089 Segment
X37089 N37089 N37090 Segment
X37090 N37090 N37091 Segment
X37091 N37091 N37092 Segment
X37092 N37092 N37093 Segment
X37093 N37093 N37094 Segment
X37094 N37094 N37095 Segment
X37095 N37095 N37096 Segment
X37096 N37096 N37097 Segment
X37097 N37097 N37098 Segment
X37098 N37098 N37099 Segment
X37099 N37099 N37100 Segment
X37100 N37100 N37101 Segment
X37101 N37101 N37102 Segment
X37102 N37102 N37103 Segment
X37103 N37103 N37104 Segment
X37104 N37104 N37105 Segment
X37105 N37105 N37106 Segment
X37106 N37106 N37107 Segment
X37107 N37107 N37108 Segment
X37108 N37108 N37109 Segment
X37109 N37109 N37110 Segment
X37110 N37110 N37111 Segment
X37111 N37111 N37112 Segment
X37112 N37112 N37113 Segment
X37113 N37113 N37114 Segment
X37114 N37114 N37115 Segment
X37115 N37115 N37116 Segment
X37116 N37116 N37117 Segment
X37117 N37117 N37118 Segment
X37118 N37118 N37119 Segment
X37119 N37119 N37120 Segment
X37120 N37120 N37121 Segment
X37121 N37121 N37122 Segment
X37122 N37122 N37123 Segment
X37123 N37123 N37124 Segment
X37124 N37124 N37125 Segment
X37125 N37125 N37126 Segment
X37126 N37126 N37127 Segment
X37127 N37127 N37128 Segment
X37128 N37128 N37129 Segment
X37129 N37129 N37130 Segment
X37130 N37130 N37131 Segment
X37131 N37131 N37132 Segment
X37132 N37132 N37133 Segment
X37133 N37133 N37134 Segment
X37134 N37134 N37135 Segment
X37135 N37135 N37136 Segment
X37136 N37136 N37137 Segment
X37137 N37137 N37138 Segment
X37138 N37138 N37139 Segment
X37139 N37139 N37140 Segment
X37140 N37140 N37141 Segment
X37141 N37141 N37142 Segment
X37142 N37142 N37143 Segment
X37143 N37143 N37144 Segment
X37144 N37144 N37145 Segment
X37145 N37145 N37146 Segment
X37146 N37146 N37147 Segment
X37147 N37147 N37148 Segment
X37148 N37148 N37149 Segment
X37149 N37149 N37150 Segment
X37150 N37150 N37151 Segment
X37151 N37151 N37152 Segment
X37152 N37152 N37153 Segment
X37153 N37153 N37154 Segment
X37154 N37154 N37155 Segment
X37155 N37155 N37156 Segment
X37156 N37156 N37157 Segment
X37157 N37157 N37158 Segment
X37158 N37158 N37159 Segment
X37159 N37159 N37160 Segment
X37160 N37160 N37161 Segment
X37161 N37161 N37162 Segment
X37162 N37162 N37163 Segment
X37163 N37163 N37164 Segment
X37164 N37164 N37165 Segment
X37165 N37165 N37166 Segment
X37166 N37166 N37167 Segment
X37167 N37167 N37168 Segment
X37168 N37168 N37169 Segment
X37169 N37169 N37170 Segment
X37170 N37170 N37171 Segment
X37171 N37171 N37172 Segment
X37172 N37172 N37173 Segment
X37173 N37173 N37174 Segment
X37174 N37174 N37175 Segment
X37175 N37175 N37176 Segment
X37176 N37176 N37177 Segment
X37177 N37177 N37178 Segment
X37178 N37178 N37179 Segment
X37179 N37179 N37180 Segment
X37180 N37180 N37181 Segment
X37181 N37181 N37182 Segment
X37182 N37182 N37183 Segment
X37183 N37183 N37184 Segment
X37184 N37184 N37185 Segment
X37185 N37185 N37186 Segment
X37186 N37186 N37187 Segment
X37187 N37187 N37188 Segment
X37188 N37188 N37189 Segment
X37189 N37189 N37190 Segment
X37190 N37190 N37191 Segment
X37191 N37191 N37192 Segment
X37192 N37192 N37193 Segment
X37193 N37193 N37194 Segment
X37194 N37194 N37195 Segment
X37195 N37195 N37196 Segment
X37196 N37196 N37197 Segment
X37197 N37197 N37198 Segment
X37198 N37198 N37199 Segment
X37199 N37199 N37200 Segment
X37200 N37200 N37201 Segment
X37201 N37201 N37202 Segment
X37202 N37202 N37203 Segment
X37203 N37203 N37204 Segment
X37204 N37204 N37205 Segment
X37205 N37205 N37206 Segment
X37206 N37206 N37207 Segment
X37207 N37207 N37208 Segment
X37208 N37208 N37209 Segment
X37209 N37209 N37210 Segment
X37210 N37210 N37211 Segment
X37211 N37211 N37212 Segment
X37212 N37212 N37213 Segment
X37213 N37213 N37214 Segment
X37214 N37214 N37215 Segment
X37215 N37215 N37216 Segment
X37216 N37216 N37217 Segment
X37217 N37217 N37218 Segment
X37218 N37218 N37219 Segment
X37219 N37219 N37220 Segment
X37220 N37220 N37221 Segment
X37221 N37221 N37222 Segment
X37222 N37222 N37223 Segment
X37223 N37223 N37224 Segment
X37224 N37224 N37225 Segment
X37225 N37225 N37226 Segment
X37226 N37226 N37227 Segment
X37227 N37227 N37228 Segment
X37228 N37228 N37229 Segment
X37229 N37229 N37230 Segment
X37230 N37230 N37231 Segment
X37231 N37231 N37232 Segment
X37232 N37232 N37233 Segment
X37233 N37233 N37234 Segment
X37234 N37234 N37235 Segment
X37235 N37235 N37236 Segment
X37236 N37236 N37237 Segment
X37237 N37237 N37238 Segment
X37238 N37238 N37239 Segment
X37239 N37239 N37240 Segment
X37240 N37240 N37241 Segment
X37241 N37241 N37242 Segment
X37242 N37242 N37243 Segment
X37243 N37243 N37244 Segment
X37244 N37244 N37245 Segment
X37245 N37245 N37246 Segment
X37246 N37246 N37247 Segment
X37247 N37247 N37248 Segment
X37248 N37248 N37249 Segment
X37249 N37249 N37250 Segment
X37250 N37250 N37251 Segment
X37251 N37251 N37252 Segment
X37252 N37252 N37253 Segment
X37253 N37253 N37254 Segment
X37254 N37254 N37255 Segment
X37255 N37255 N37256 Segment
X37256 N37256 N37257 Segment
X37257 N37257 N37258 Segment
X37258 N37258 N37259 Segment
X37259 N37259 N37260 Segment
X37260 N37260 N37261 Segment
X37261 N37261 N37262 Segment
X37262 N37262 N37263 Segment
X37263 N37263 N37264 Segment
X37264 N37264 N37265 Segment
X37265 N37265 N37266 Segment
X37266 N37266 N37267 Segment
X37267 N37267 N37268 Segment
X37268 N37268 N37269 Segment
X37269 N37269 N37270 Segment
X37270 N37270 N37271 Segment
X37271 N37271 N37272 Segment
X37272 N37272 N37273 Segment
X37273 N37273 N37274 Segment
X37274 N37274 N37275 Segment
X37275 N37275 N37276 Segment
X37276 N37276 N37277 Segment
X37277 N37277 N37278 Segment
X37278 N37278 N37279 Segment
X37279 N37279 N37280 Segment
X37280 N37280 N37281 Segment
X37281 N37281 N37282 Segment
X37282 N37282 N37283 Segment
X37283 N37283 N37284 Segment
X37284 N37284 N37285 Segment
X37285 N37285 N37286 Segment
X37286 N37286 N37287 Segment
X37287 N37287 N37288 Segment
X37288 N37288 N37289 Segment
X37289 N37289 N37290 Segment
X37290 N37290 N37291 Segment
X37291 N37291 N37292 Segment
X37292 N37292 N37293 Segment
X37293 N37293 N37294 Segment
X37294 N37294 N37295 Segment
X37295 N37295 N37296 Segment
X37296 N37296 N37297 Segment
X37297 N37297 N37298 Segment
X37298 N37298 N37299 Segment
X37299 N37299 N37300 Segment
X37300 N37300 N37301 Segment
X37301 N37301 N37302 Segment
X37302 N37302 N37303 Segment
X37303 N37303 N37304 Segment
X37304 N37304 N37305 Segment
X37305 N37305 N37306 Segment
X37306 N37306 N37307 Segment
X37307 N37307 N37308 Segment
X37308 N37308 N37309 Segment
X37309 N37309 N37310 Segment
X37310 N37310 N37311 Segment
X37311 N37311 N37312 Segment
X37312 N37312 N37313 Segment
X37313 N37313 N37314 Segment
X37314 N37314 N37315 Segment
X37315 N37315 N37316 Segment
X37316 N37316 N37317 Segment
X37317 N37317 N37318 Segment
X37318 N37318 N37319 Segment
X37319 N37319 N37320 Segment
X37320 N37320 N37321 Segment
X37321 N37321 N37322 Segment
X37322 N37322 N37323 Segment
X37323 N37323 N37324 Segment
X37324 N37324 N37325 Segment
X37325 N37325 N37326 Segment
X37326 N37326 N37327 Segment
X37327 N37327 N37328 Segment
X37328 N37328 N37329 Segment
X37329 N37329 N37330 Segment
X37330 N37330 N37331 Segment
X37331 N37331 N37332 Segment
X37332 N37332 N37333 Segment
X37333 N37333 N37334 Segment
X37334 N37334 N37335 Segment
X37335 N37335 N37336 Segment
X37336 N37336 N37337 Segment
X37337 N37337 N37338 Segment
X37338 N37338 N37339 Segment
X37339 N37339 N37340 Segment
X37340 N37340 N37341 Segment
X37341 N37341 N37342 Segment
X37342 N37342 N37343 Segment
X37343 N37343 N37344 Segment
X37344 N37344 N37345 Segment
X37345 N37345 N37346 Segment
X37346 N37346 N37347 Segment
X37347 N37347 N37348 Segment
X37348 N37348 N37349 Segment
X37349 N37349 N37350 Segment
X37350 N37350 N37351 Segment
X37351 N37351 N37352 Segment
X37352 N37352 N37353 Segment
X37353 N37353 N37354 Segment
X37354 N37354 N37355 Segment
X37355 N37355 N37356 Segment
X37356 N37356 N37357 Segment
X37357 N37357 N37358 Segment
X37358 N37358 N37359 Segment
X37359 N37359 N37360 Segment
X37360 N37360 N37361 Segment
X37361 N37361 N37362 Segment
X37362 N37362 N37363 Segment
X37363 N37363 N37364 Segment
X37364 N37364 N37365 Segment
X37365 N37365 N37366 Segment
X37366 N37366 N37367 Segment
X37367 N37367 N37368 Segment
X37368 N37368 N37369 Segment
X37369 N37369 N37370 Segment
X37370 N37370 N37371 Segment
X37371 N37371 N37372 Segment
X37372 N37372 N37373 Segment
X37373 N37373 N37374 Segment
X37374 N37374 N37375 Segment
X37375 N37375 N37376 Segment
X37376 N37376 N37377 Segment
X37377 N37377 N37378 Segment
X37378 N37378 N37379 Segment
X37379 N37379 N37380 Segment
X37380 N37380 N37381 Segment
X37381 N37381 N37382 Segment
X37382 N37382 N37383 Segment
X37383 N37383 N37384 Segment
X37384 N37384 N37385 Segment
X37385 N37385 N37386 Segment
X37386 N37386 N37387 Segment
X37387 N37387 N37388 Segment
X37388 N37388 N37389 Segment
X37389 N37389 N37390 Segment
X37390 N37390 N37391 Segment
X37391 N37391 N37392 Segment
X37392 N37392 N37393 Segment
X37393 N37393 N37394 Segment
X37394 N37394 N37395 Segment
X37395 N37395 N37396 Segment
X37396 N37396 N37397 Segment
X37397 N37397 N37398 Segment
X37398 N37398 N37399 Segment
X37399 N37399 N37400 Segment
X37400 N37400 N37401 Segment
X37401 N37401 N37402 Segment
X37402 N37402 N37403 Segment
X37403 N37403 N37404 Segment
X37404 N37404 N37405 Segment
X37405 N37405 N37406 Segment
X37406 N37406 N37407 Segment
X37407 N37407 N37408 Segment
X37408 N37408 N37409 Segment
X37409 N37409 N37410 Segment
X37410 N37410 N37411 Segment
X37411 N37411 N37412 Segment
X37412 N37412 N37413 Segment
X37413 N37413 N37414 Segment
X37414 N37414 N37415 Segment
X37415 N37415 N37416 Segment
X37416 N37416 N37417 Segment
X37417 N37417 N37418 Segment
X37418 N37418 N37419 Segment
X37419 N37419 N37420 Segment
X37420 N37420 N37421 Segment
X37421 N37421 N37422 Segment
X37422 N37422 N37423 Segment
X37423 N37423 N37424 Segment
X37424 N37424 N37425 Segment
X37425 N37425 N37426 Segment
X37426 N37426 N37427 Segment
X37427 N37427 N37428 Segment
X37428 N37428 N37429 Segment
X37429 N37429 N37430 Segment
X37430 N37430 N37431 Segment
X37431 N37431 N37432 Segment
X37432 N37432 N37433 Segment
X37433 N37433 N37434 Segment
X37434 N37434 N37435 Segment
X37435 N37435 N37436 Segment
X37436 N37436 N37437 Segment
X37437 N37437 N37438 Segment
X37438 N37438 N37439 Segment
X37439 N37439 N37440 Segment
X37440 N37440 N37441 Segment
X37441 N37441 N37442 Segment
X37442 N37442 N37443 Segment
X37443 N37443 N37444 Segment
X37444 N37444 N37445 Segment
X37445 N37445 N37446 Segment
X37446 N37446 N37447 Segment
X37447 N37447 N37448 Segment
X37448 N37448 N37449 Segment
X37449 N37449 N37450 Segment
X37450 N37450 N37451 Segment
X37451 N37451 N37452 Segment
X37452 N37452 N37453 Segment
X37453 N37453 N37454 Segment
X37454 N37454 N37455 Segment
X37455 N37455 N37456 Segment
X37456 N37456 N37457 Segment
X37457 N37457 N37458 Segment
X37458 N37458 N37459 Segment
X37459 N37459 N37460 Segment
X37460 N37460 N37461 Segment
X37461 N37461 N37462 Segment
X37462 N37462 N37463 Segment
X37463 N37463 N37464 Segment
X37464 N37464 N37465 Segment
X37465 N37465 N37466 Segment
X37466 N37466 N37467 Segment
X37467 N37467 N37468 Segment
X37468 N37468 N37469 Segment
X37469 N37469 N37470 Segment
X37470 N37470 N37471 Segment
X37471 N37471 N37472 Segment
X37472 N37472 N37473 Segment
X37473 N37473 N37474 Segment
X37474 N37474 N37475 Segment
X37475 N37475 N37476 Segment
X37476 N37476 N37477 Segment
X37477 N37477 N37478 Segment
X37478 N37478 N37479 Segment
X37479 N37479 N37480 Segment
X37480 N37480 N37481 Segment
X37481 N37481 N37482 Segment
X37482 N37482 N37483 Segment
X37483 N37483 N37484 Segment
X37484 N37484 N37485 Segment
X37485 N37485 N37486 Segment
X37486 N37486 N37487 Segment
X37487 N37487 N37488 Segment
X37488 N37488 N37489 Segment
X37489 N37489 N37490 Segment
X37490 N37490 N37491 Segment
X37491 N37491 N37492 Segment
X37492 N37492 N37493 Segment
X37493 N37493 N37494 Segment
X37494 N37494 N37495 Segment
X37495 N37495 N37496 Segment
X37496 N37496 N37497 Segment
X37497 N37497 N37498 Segment
X37498 N37498 N37499 Segment
X37499 N37499 N37500 Segment
X37500 N37500 N37501 Segment
X37501 N37501 N37502 Segment
X37502 N37502 N37503 Segment
X37503 N37503 N37504 Segment
X37504 N37504 N37505 Segment
X37505 N37505 N37506 Segment
X37506 N37506 N37507 Segment
X37507 N37507 N37508 Segment
X37508 N37508 N37509 Segment
X37509 N37509 N37510 Segment
X37510 N37510 N37511 Segment
X37511 N37511 N37512 Segment
X37512 N37512 N37513 Segment
X37513 N37513 N37514 Segment
X37514 N37514 N37515 Segment
X37515 N37515 N37516 Segment
X37516 N37516 N37517 Segment
X37517 N37517 N37518 Segment
X37518 N37518 N37519 Segment
X37519 N37519 N37520 Segment
X37520 N37520 N37521 Segment
X37521 N37521 N37522 Segment
X37522 N37522 N37523 Segment
X37523 N37523 N37524 Segment
X37524 N37524 N37525 Segment
X37525 N37525 N37526 Segment
X37526 N37526 N37527 Segment
X37527 N37527 N37528 Segment
X37528 N37528 N37529 Segment
X37529 N37529 N37530 Segment
X37530 N37530 N37531 Segment
X37531 N37531 N37532 Segment
X37532 N37532 N37533 Segment
X37533 N37533 N37534 Segment
X37534 N37534 N37535 Segment
X37535 N37535 N37536 Segment
X37536 N37536 N37537 Segment
X37537 N37537 N37538 Segment
X37538 N37538 N37539 Segment
X37539 N37539 N37540 Segment
X37540 N37540 N37541 Segment
X37541 N37541 N37542 Segment
X37542 N37542 N37543 Segment
X37543 N37543 N37544 Segment
X37544 N37544 N37545 Segment
X37545 N37545 N37546 Segment
X37546 N37546 N37547 Segment
X37547 N37547 N37548 Segment
X37548 N37548 Vout Segment

* Source and load
V1 Vsource 0 PULSE(0 10 0 5.0e-13 5.0e-13 5n)
Rsource Vsource Vin 50
Rload Vout 0 121.3

* Simulation command
.tran 20n
.end
